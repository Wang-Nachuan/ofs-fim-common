// Copyright 2021 Intel Corporation
// SPDX-License-Identifier: MIT

`include "fim_gram_sdp.v"
`include "fim_ram_1r1w.sv"
`include "bfifo.sv"
`include "pfa_master.sv"
`include "pfa_master_tb.sv"
