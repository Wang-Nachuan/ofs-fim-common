// Copyright (C) 2023 Intel Corporation
// SPDX-License-Identifier: MIT

`include "svt_axi.uvm.pkg"
`include "uvm_pkg.sv"
`include "sequence_lib.svh"
`include "test_package.sv"

`ifdef TB_CONFIG_1
`define NUM_PORT 16;
localparam LOCAL_NUM_RTABLE_ENTRIES = 16;
 `ifdef INVALID_PF_VF  //{
   localparam pf_vf_mux_pkg::t_pfvf_rtable_entry LOCAL_PFVF_ROUTING_TABLE[LOCAL_NUM_RTABLE_ENTRIES] = '{
            '{ pfvf_port:0 , pf:0 , vf:0 , vf_active:0  },         // PF0 to PF7
            '{ pfvf_port:1 , pf:1 , vf:0 , vf_active:0  },
            '{ pfvf_port:2 , pf:2 , vf:0 , vf_active:0  },
            '{ pfvf_port:3 , pf:3 , vf:0 , vf_active:0  },
            '{ pfvf_port:4 , pf:4 , vf:0 , vf_active:0  },
            '{ pfvf_port:5 , pf:5 , vf:0 , vf_active:0  },
            '{ pfvf_port:6 , pf:6 , vf:0 , vf_active:0  },
            '{ pfvf_port:7 , pf:7 , vf:0 , vf_active:0  },
            '{ pfvf_port:8 , pf:0 , vf:3 , vf_active:1  },        // PF0-VF0 to PF7-VF0 
            '{ pfvf_port:9 , pf:1 , vf:3 , vf_active:1  },
            '{ pfvf_port:10 , pf:2 , vf:3 , vf_active:1  },
            '{ pfvf_port:11 , pf:3 , vf:3 , vf_active:1  },
            '{ pfvf_port:12 , pf:4 , vf:3 , vf_active:1  },
            '{ pfvf_port:13 , pf:5 , vf:3 , vf_active:1  },
            '{ pfvf_port:14 , pf:6 , vf:3 , vf_active:1  },
            '{ pfvf_port:15 , pf:7 , vf:3 , vf_active:1  }
          };
  `else
    localparam pf_vf_mux_pkg::t_pfvf_rtable_entry LOCAL_PFVF_ROUTING_TABLE[LOCAL_NUM_RTABLE_ENTRIES] = '{
            '{ pfvf_port:0 , pf:0 , vf:0 , vf_active:0  },         // PF0 to PF7
            '{ pfvf_port:1 , pf:1 , vf:0 , vf_active:0  },
            '{ pfvf_port:2 , pf:2 , vf:0 , vf_active:0  },
            '{ pfvf_port:3 , pf:3 , vf:0 , vf_active:0  },
            '{ pfvf_port:4 , pf:4 , vf:0 , vf_active:0  },
            '{ pfvf_port:5 , pf:5 , vf:0 , vf_active:0  },
            '{ pfvf_port:6 , pf:6 , vf:0 , vf_active:0  },
            '{ pfvf_port:7 , pf:7 , vf:0 , vf_active:0  },
            '{ pfvf_port:8 , pf:0 , vf:0 , vf_active:1  },        // PF0-VF0 to PF7-VF0 
            '{ pfvf_port:9 , pf:1 , vf:0 , vf_active:1  },
            '{ pfvf_port:10 , pf:2 , vf:0 , vf_active:1  },
            '{ pfvf_port:11 , pf:3 , vf:0 , vf_active:1  },
            '{ pfvf_port:12 , pf:4 , vf:0 , vf_active:1  },
            '{ pfvf_port:13 , pf:5 , vf:0 , vf_active:1  },
            '{ pfvf_port:14 , pf:6 , vf:0 , vf_active:1  },
            '{ pfvf_port:15 , pf:7 , vf:0 , vf_active:1  }
          };
  `endif  //}
`elsif TB_CONFIG_2
`define NUM_PORT 24;
localparam LOCAL_NUM_RTABLE_ENTRIES = 24;
localparam pf_vf_mux_pkg::t_pfvf_rtable_entry LOCAL_PFVF_ROUTING_TABLE[LOCAL_NUM_RTABLE_ENTRIES] = '{
          '{ pfvf_port:0  , pf:0 , vf:0    , vf_active:0  },      // PF0 to PF7
          '{ pfvf_port:1  , pf:1 , vf:0    , vf_active:0  },
          '{ pfvf_port:2  , pf:2 , vf:0    , vf_active:0  },
          '{ pfvf_port:3  , pf:3 , vf:0    , vf_active:0  },
          '{ pfvf_port:4  , pf:4 , vf:0    , vf_active:0  },
          '{ pfvf_port:5  , pf:5 , vf:0    , vf_active:0  },
          '{ pfvf_port:6  , pf:6 , vf:0    , vf_active:0  },
          '{ pfvf_port:7  , pf:7 , vf:0    , vf_active:0  },
          '{ pfvf_port:8  , pf:0 , vf:0    , vf_active:1  },     // PF0-VF0 to PF7-VF0
          '{ pfvf_port:9  , pf:1 , vf:0    , vf_active:1  }, 
          '{ pfvf_port:10 , pf:2 , vf:0    , vf_active:1  },
          '{ pfvf_port:11 , pf:3 , vf:0    , vf_active:1  },
          '{ pfvf_port:12 , pf:4 , vf:0    , vf_active:1  },
          '{ pfvf_port:13 , pf:5 , vf:0    , vf_active:1  },
          '{ pfvf_port:14 , pf:6 , vf:0    , vf_active:1  },
          '{ pfvf_port:15 , pf:7 , vf:0    , vf_active:1  },
          '{ pfvf_port:16 , pf:0 , vf:2047 , vf_active:1  },     // PF0-VF2047 to PF7-VF2047
          '{ pfvf_port:17 , pf:1 , vf:2047 , vf_active:1  },
          '{ pfvf_port:18 , pf:2 , vf:2047 , vf_active:1  },
          '{ pfvf_port:19 , pf:3 , vf:2047 , vf_active:1  },
          '{ pfvf_port:20 , pf:4 , vf:2047 , vf_active:1  },
          '{ pfvf_port:21 , pf:5 , vf:2047 , vf_active:1  },
          '{ pfvf_port:22 , pf:6 , vf:2047 , vf_active:1  },
          '{ pfvf_port:23 , pf:7 , vf:2047 , vf_active:1  }
        };
`elsif TB_CONFIG_3
`define NUM_PORT 32;
localparam LOCAL_NUM_RTABLE_ENTRIES = 32;
localparam pf_vf_mux_pkg::t_pfvf_rtable_entry LOCAL_PFVF_ROUTING_TABLE[LOCAL_NUM_RTABLE_ENTRIES] = '{
          '{ pfvf_port:0  , pf:0 , vf:0    , vf_active:0  },      // PF0 to PF7
          '{ pfvf_port:1  , pf:1 , vf:0    , vf_active:0  },
          '{ pfvf_port:2  , pf:2 , vf:0    , vf_active:0  },
          '{ pfvf_port:3  , pf:3 , vf:0    , vf_active:0  },
          '{ pfvf_port:4  , pf:4 , vf:0    , vf_active:0  },
          '{ pfvf_port:5  , pf:5 , vf:0    , vf_active:0  },
          '{ pfvf_port:6  , pf:6 , vf:0    , vf_active:0  },
          '{ pfvf_port:7  , pf:7 , vf:0    , vf_active:0  },
          '{ pfvf_port:8  , pf:0 , vf:0    , vf_active:1  },     // PF0-VF0 to PF7-VF0
          '{ pfvf_port:9  , pf:1 , vf:0    , vf_active:1  }, 
          '{ pfvf_port:10 , pf:2 , vf:0    , vf_active:1  },
          '{ pfvf_port:11 , pf:3 , vf:0    , vf_active:1  },
          '{ pfvf_port:12 , pf:4 , vf:0    , vf_active:1  },
          '{ pfvf_port:13 , pf:5 , vf:0    , vf_active:1  },
          '{ pfvf_port:14 , pf:6 , vf:0    , vf_active:1  },
          '{ pfvf_port:15 , pf:7 , vf:0    , vf_active:1  },
          '{ pfvf_port:16 , pf:0 , vf:2047 , vf_active:1  },     // PF0-VF2047 to PF7-VF2047
          '{ pfvf_port:17 , pf:1 , vf:2047 , vf_active:1  },
          '{ pfvf_port:18 , pf:2 , vf:2047 , vf_active:1  },
          '{ pfvf_port:19 , pf:3 , vf:2047 , vf_active:1  },
          '{ pfvf_port:20 , pf:4 , vf:2047 , vf_active:1  },
          '{ pfvf_port:21 , pf:5 , vf:2047 , vf_active:1  },
          '{ pfvf_port:22 , pf:6 , vf:2047 , vf_active:1  },
          '{ pfvf_port:23 , pf:7 , vf:2047 , vf_active:1  },
          '{ pfvf_port:24 , pf:0 , vf:`RANDOM_VF   , vf_active:1  },
          '{ pfvf_port:25 , pf:1 , vf:`RANDOM_VF   , vf_active:1  },
          '{ pfvf_port:26 , pf:2 , vf:`RANDOM_VF   , vf_active:1  },
          '{ pfvf_port:27 , pf:3 , vf:`RANDOM_VF   , vf_active:1  },
          '{ pfvf_port:28 , pf:4 , vf:`RANDOM_VF   , vf_active:1  },
          '{ pfvf_port:29 , pf:5 , vf:`RANDOM_VF   , vf_active:1  },
          '{ pfvf_port:30 , pf:6 , vf:`RANDOM_VF   , vf_active:1  },
          '{ pfvf_port:31 , pf:7 , vf:`RANDOM_VF   , vf_active:1  }
        };
`elsif TB_CONFIG_4
`define NUM_PORT 2048;
localparam LOCAL_NUM_RTABLE_ENTRIES = 2048;
localparam pf_vf_mux_pkg::t_pfvf_rtable_entry [LOCAL_NUM_RTABLE_ENTRIES-1:0] LOCAL_PFVF_ROUTING_TABLE = '{
'{ pfvf_port:0  , pf:0 , vf:0    , vf_active:1  },      
'{ pfvf_port:1  , pf:0 , vf:1    , vf_active:1  },      
'{ pfvf_port:2  , pf:0 , vf:2    , vf_active:1  },      
'{ pfvf_port:3  , pf:0 , vf:3    , vf_active:1  },      
'{ pfvf_port:4  , pf:0 , vf:4    , vf_active:1  },      
'{ pfvf_port:5  , pf:0 , vf:5    , vf_active:1  },      
'{ pfvf_port:6  , pf:0 , vf:6    , vf_active:1  },      
'{ pfvf_port:7  , pf:0 , vf:7    , vf_active:1  },      
'{ pfvf_port:8  , pf:0 , vf:8    , vf_active:1  },      
'{ pfvf_port:9  , pf:0 , vf:9    , vf_active:1  },      
'{ pfvf_port:10  , pf:0 , vf:10    , vf_active:1  },      
'{ pfvf_port:11  , pf:0 , vf:11    , vf_active:1  },      
'{ pfvf_port:12  , pf:0 , vf:12    , vf_active:1  },      
'{ pfvf_port:13  , pf:0 , vf:13    , vf_active:1  },      
'{ pfvf_port:14  , pf:0 , vf:14    , vf_active:1  },      
'{ pfvf_port:15  , pf:0 , vf:15    , vf_active:1  },      
'{ pfvf_port:16  , pf:0 , vf:16    , vf_active:1  },      
'{ pfvf_port:17  , pf:0 , vf:17    , vf_active:1  },      
'{ pfvf_port:18  , pf:0 , vf:18    , vf_active:1  },      
'{ pfvf_port:19  , pf:0 , vf:19    , vf_active:1  },      
'{ pfvf_port:20  , pf:0 , vf:20    , vf_active:1  },      
'{ pfvf_port:21  , pf:0 , vf:21    , vf_active:1  },      
'{ pfvf_port:22  , pf:0 , vf:22    , vf_active:1  },      
'{ pfvf_port:23  , pf:0 , vf:23    , vf_active:1  },      
'{ pfvf_port:24  , pf:0 , vf:24    , vf_active:1  },      
'{ pfvf_port:25  , pf:0 , vf:25    , vf_active:1  },      
'{ pfvf_port:26  , pf:0 , vf:26    , vf_active:1  },      
'{ pfvf_port:27  , pf:0 , vf:27    , vf_active:1  },      
'{ pfvf_port:28  , pf:0 , vf:28    , vf_active:1  },      
'{ pfvf_port:29  , pf:0 , vf:29    , vf_active:1  },      
'{ pfvf_port:30  , pf:0 , vf:30    , vf_active:1  },      
'{ pfvf_port:31  , pf:0 , vf:31    , vf_active:1  },      
'{ pfvf_port:32  , pf:0 , vf:32    , vf_active:1  },      
'{ pfvf_port:33  , pf:0 , vf:33    , vf_active:1  },      
'{ pfvf_port:34  , pf:0 , vf:34    , vf_active:1  },      
'{ pfvf_port:35  , pf:0 , vf:35    , vf_active:1  },      
'{ pfvf_port:36  , pf:0 , vf:36    , vf_active:1  },      
'{ pfvf_port:37  , pf:0 , vf:37    , vf_active:1  },      
'{ pfvf_port:38  , pf:0 , vf:38    , vf_active:1  },      
'{ pfvf_port:39  , pf:0 , vf:39    , vf_active:1  },      
'{ pfvf_port:40  , pf:0 , vf:40    , vf_active:1  },      
'{ pfvf_port:41  , pf:0 , vf:41    , vf_active:1  },      
'{ pfvf_port:42  , pf:0 , vf:42    , vf_active:1  },      
'{ pfvf_port:43  , pf:0 , vf:43    , vf_active:1  },      
'{ pfvf_port:44  , pf:0 , vf:44    , vf_active:1  },      
'{ pfvf_port:45  , pf:0 , vf:45    , vf_active:1  },      
'{ pfvf_port:46  , pf:0 , vf:46    , vf_active:1  },      
'{ pfvf_port:47  , pf:0 , vf:47    , vf_active:1  },      
'{ pfvf_port:48  , pf:0 , vf:48    , vf_active:1  },      
'{ pfvf_port:49  , pf:0 , vf:49    , vf_active:1  },      
'{ pfvf_port:50  , pf:0 , vf:50    , vf_active:1  },      
'{ pfvf_port:51  , pf:0 , vf:51    , vf_active:1  },      
'{ pfvf_port:52  , pf:0 , vf:52    , vf_active:1  },      
'{ pfvf_port:53  , pf:0 , vf:53    , vf_active:1  },      
'{ pfvf_port:54  , pf:0 , vf:54    , vf_active:1  },      
'{ pfvf_port:55  , pf:0 , vf:55    , vf_active:1  },      
'{ pfvf_port:56  , pf:0 , vf:56    , vf_active:1  },      
'{ pfvf_port:57  , pf:0 , vf:57    , vf_active:1  },      
'{ pfvf_port:58  , pf:0 , vf:58    , vf_active:1  },      
'{ pfvf_port:59  , pf:0 , vf:59    , vf_active:1  },      
'{ pfvf_port:60  , pf:0 , vf:60    , vf_active:1  },      
'{ pfvf_port:61  , pf:0 , vf:61    , vf_active:1  },      
'{ pfvf_port:62  , pf:0 , vf:62    , vf_active:1  },      
'{ pfvf_port:63  , pf:0 , vf:63    , vf_active:1  },      
'{ pfvf_port:64  , pf:0 , vf:64    , vf_active:1  },      
'{ pfvf_port:65  , pf:0 , vf:65    , vf_active:1  },      
'{ pfvf_port:66  , pf:0 , vf:66    , vf_active:1  },      
'{ pfvf_port:67  , pf:0 , vf:67    , vf_active:1  },      
'{ pfvf_port:68  , pf:0 , vf:68    , vf_active:1  },      
'{ pfvf_port:69  , pf:0 , vf:69    , vf_active:1  },      
'{ pfvf_port:70  , pf:0 , vf:70    , vf_active:1  },      
'{ pfvf_port:71  , pf:0 , vf:71    , vf_active:1  },      
'{ pfvf_port:72  , pf:0 , vf:72    , vf_active:1  },      
'{ pfvf_port:73  , pf:0 , vf:73    , vf_active:1  },      
'{ pfvf_port:74  , pf:0 , vf:74    , vf_active:1  },      
'{ pfvf_port:75  , pf:0 , vf:75    , vf_active:1  },      
'{ pfvf_port:76  , pf:0 , vf:76    , vf_active:1  },      
'{ pfvf_port:77  , pf:0 , vf:77    , vf_active:1  },      
'{ pfvf_port:78  , pf:0 , vf:78    , vf_active:1  },      
'{ pfvf_port:79  , pf:0 , vf:79    , vf_active:1  },      
'{ pfvf_port:80  , pf:0 , vf:80    , vf_active:1  },      
'{ pfvf_port:81  , pf:0 , vf:81    , vf_active:1  },      
'{ pfvf_port:82  , pf:0 , vf:82    , vf_active:1  },      
'{ pfvf_port:83  , pf:0 , vf:83    , vf_active:1  },      
'{ pfvf_port:84  , pf:0 , vf:84    , vf_active:1  },      
'{ pfvf_port:85  , pf:0 , vf:85    , vf_active:1  },      
'{ pfvf_port:86  , pf:0 , vf:86    , vf_active:1  },      
'{ pfvf_port:87  , pf:0 , vf:87    , vf_active:1  },      
'{ pfvf_port:88  , pf:0 , vf:88    , vf_active:1  },      
'{ pfvf_port:89  , pf:0 , vf:89    , vf_active:1  },      
'{ pfvf_port:90  , pf:0 , vf:90    , vf_active:1  },      
'{ pfvf_port:91  , pf:0 , vf:91    , vf_active:1  },      
'{ pfvf_port:92  , pf:0 , vf:92    , vf_active:1  },      
'{ pfvf_port:93  , pf:0 , vf:93    , vf_active:1  },      
'{ pfvf_port:94  , pf:0 , vf:94    , vf_active:1  },      
'{ pfvf_port:95  , pf:0 , vf:95    , vf_active:1  },      
'{ pfvf_port:96  , pf:0 , vf:96    , vf_active:1  },      
'{ pfvf_port:97  , pf:0 , vf:97    , vf_active:1  },      
'{ pfvf_port:98  , pf:0 , vf:98    , vf_active:1  },      
'{ pfvf_port:99  , pf:0 , vf:99    , vf_active:1  },      
'{ pfvf_port:100  , pf:0 , vf:100    , vf_active:1  },      
'{ pfvf_port:101  , pf:0 , vf:101    , vf_active:1  },      
'{ pfvf_port:102  , pf:0 , vf:102    , vf_active:1  },      
'{ pfvf_port:103  , pf:0 , vf:103    , vf_active:1  },      
'{ pfvf_port:104  , pf:0 , vf:104    , vf_active:1  },      
'{ pfvf_port:105  , pf:0 , vf:105    , vf_active:1  },      
'{ pfvf_port:106  , pf:0 , vf:106    , vf_active:1  },      
'{ pfvf_port:107  , pf:0 , vf:107    , vf_active:1  },      
'{ pfvf_port:108  , pf:0 , vf:108    , vf_active:1  },      
'{ pfvf_port:109  , pf:0 , vf:109    , vf_active:1  },      
'{ pfvf_port:110  , pf:0 , vf:110    , vf_active:1  },      
'{ pfvf_port:111  , pf:0 , vf:111    , vf_active:1  },      
'{ pfvf_port:112  , pf:0 , vf:112    , vf_active:1  },      
'{ pfvf_port:113  , pf:0 , vf:113    , vf_active:1  },      
'{ pfvf_port:114  , pf:0 , vf:114    , vf_active:1  },      
'{ pfvf_port:115  , pf:0 , vf:115    , vf_active:1  },      
'{ pfvf_port:116  , pf:0 , vf:116    , vf_active:1  },      
'{ pfvf_port:117  , pf:0 , vf:117    , vf_active:1  },      
'{ pfvf_port:118  , pf:0 , vf:118    , vf_active:1  },      
'{ pfvf_port:119  , pf:0 , vf:119    , vf_active:1  },      
'{ pfvf_port:120  , pf:0 , vf:120    , vf_active:1  },      
'{ pfvf_port:121  , pf:0 , vf:121    , vf_active:1  },      
'{ pfvf_port:122  , pf:0 , vf:122    , vf_active:1  },      
'{ pfvf_port:123  , pf:0 , vf:123    , vf_active:1  },      
'{ pfvf_port:124  , pf:0 , vf:124    , vf_active:1  },      
'{ pfvf_port:125  , pf:0 , vf:125    , vf_active:1  },      
'{ pfvf_port:126  , pf:0 , vf:126    , vf_active:1  },      
'{ pfvf_port:127  , pf:0 , vf:127    , vf_active:1  },      
'{ pfvf_port:128  , pf:0 , vf:128    , vf_active:1  },      
'{ pfvf_port:129  , pf:0 , vf:129    , vf_active:1  },      
'{ pfvf_port:130  , pf:0 , vf:130    , vf_active:1  },      
'{ pfvf_port:131  , pf:0 , vf:131    , vf_active:1  },      
'{ pfvf_port:132  , pf:0 , vf:132    , vf_active:1  },      
'{ pfvf_port:133  , pf:0 , vf:133    , vf_active:1  },      
'{ pfvf_port:134  , pf:0 , vf:134    , vf_active:1  },      
'{ pfvf_port:135  , pf:0 , vf:135    , vf_active:1  },      
'{ pfvf_port:136  , pf:0 , vf:136    , vf_active:1  },      
'{ pfvf_port:137  , pf:0 , vf:137    , vf_active:1  },      
'{ pfvf_port:138  , pf:0 , vf:138    , vf_active:1  },      
'{ pfvf_port:139  , pf:0 , vf:139    , vf_active:1  },      
'{ pfvf_port:140  , pf:0 , vf:140    , vf_active:1  },      
'{ pfvf_port:141  , pf:0 , vf:141    , vf_active:1  },      
'{ pfvf_port:142  , pf:0 , vf:142    , vf_active:1  },      
'{ pfvf_port:143  , pf:0 , vf:143    , vf_active:1  },      
'{ pfvf_port:144  , pf:0 , vf:144    , vf_active:1  },      
'{ pfvf_port:145  , pf:0 , vf:145    , vf_active:1  },      
'{ pfvf_port:146  , pf:0 , vf:146    , vf_active:1  },      
'{ pfvf_port:147  , pf:0 , vf:147    , vf_active:1  },      
'{ pfvf_port:148  , pf:0 , vf:148    , vf_active:1  },      
'{ pfvf_port:149  , pf:0 , vf:149    , vf_active:1  },      
'{ pfvf_port:150  , pf:0 , vf:150    , vf_active:1  },      
'{ pfvf_port:151  , pf:0 , vf:151    , vf_active:1  },      
'{ pfvf_port:152  , pf:0 , vf:152    , vf_active:1  },      
'{ pfvf_port:153  , pf:0 , vf:153    , vf_active:1  },      
'{ pfvf_port:154  , pf:0 , vf:154    , vf_active:1  },      
'{ pfvf_port:155  , pf:0 , vf:155    , vf_active:1  },      
'{ pfvf_port:156  , pf:0 , vf:156    , vf_active:1  },      
'{ pfvf_port:157  , pf:0 , vf:157    , vf_active:1  },      
'{ pfvf_port:158  , pf:0 , vf:158    , vf_active:1  },      
'{ pfvf_port:159  , pf:0 , vf:159    , vf_active:1  },      
'{ pfvf_port:160  , pf:0 , vf:160    , vf_active:1  },      
'{ pfvf_port:161  , pf:0 , vf:161    , vf_active:1  },      
'{ pfvf_port:162  , pf:0 , vf:162    , vf_active:1  },      
'{ pfvf_port:163  , pf:0 , vf:163    , vf_active:1  },      
'{ pfvf_port:164  , pf:0 , vf:164    , vf_active:1  },      
'{ pfvf_port:165  , pf:0 , vf:165    , vf_active:1  },      
'{ pfvf_port:166  , pf:0 , vf:166    , vf_active:1  },      
'{ pfvf_port:167  , pf:0 , vf:167    , vf_active:1  },      
'{ pfvf_port:168  , pf:0 , vf:168    , vf_active:1  },      
'{ pfvf_port:169  , pf:0 , vf:169    , vf_active:1  },      
'{ pfvf_port:170  , pf:0 , vf:170    , vf_active:1  },      
'{ pfvf_port:171  , pf:0 , vf:171    , vf_active:1  },      
'{ pfvf_port:172  , pf:0 , vf:172    , vf_active:1  },      
'{ pfvf_port:173  , pf:0 , vf:173    , vf_active:1  },      
'{ pfvf_port:174  , pf:0 , vf:174    , vf_active:1  },      
'{ pfvf_port:175  , pf:0 , vf:175    , vf_active:1  },      
'{ pfvf_port:176  , pf:0 , vf:176    , vf_active:1  },      
'{ pfvf_port:177  , pf:0 , vf:177    , vf_active:1  },      
'{ pfvf_port:178  , pf:0 , vf:178    , vf_active:1  },      
'{ pfvf_port:179  , pf:0 , vf:179    , vf_active:1  },      
'{ pfvf_port:180  , pf:0 , vf:180    , vf_active:1  },      
'{ pfvf_port:181  , pf:0 , vf:181    , vf_active:1  },      
'{ pfvf_port:182  , pf:0 , vf:182    , vf_active:1  },      
'{ pfvf_port:183  , pf:0 , vf:183    , vf_active:1  },      
'{ pfvf_port:184  , pf:0 , vf:184    , vf_active:1  },      
'{ pfvf_port:185  , pf:0 , vf:185    , vf_active:1  },      
'{ pfvf_port:186  , pf:0 , vf:186    , vf_active:1  },      
'{ pfvf_port:187  , pf:0 , vf:187    , vf_active:1  },      
'{ pfvf_port:188  , pf:0 , vf:188    , vf_active:1  },      
'{ pfvf_port:189  , pf:0 , vf:189    , vf_active:1  },      
'{ pfvf_port:190  , pf:0 , vf:190    , vf_active:1  },      
'{ pfvf_port:191  , pf:0 , vf:191    , vf_active:1  },      
'{ pfvf_port:192  , pf:0 , vf:192    , vf_active:1  },      
'{ pfvf_port:193  , pf:0 , vf:193    , vf_active:1  },      
'{ pfvf_port:194  , pf:0 , vf:194    , vf_active:1  },      
'{ pfvf_port:195  , pf:0 , vf:195    , vf_active:1  },      
'{ pfvf_port:196  , pf:0 , vf:196    , vf_active:1  },      
'{ pfvf_port:197  , pf:0 , vf:197    , vf_active:1  },      
'{ pfvf_port:198  , pf:0 , vf:198    , vf_active:1  },      
'{ pfvf_port:199  , pf:0 , vf:199    , vf_active:1  },      
'{ pfvf_port:200  , pf:0 , vf:200    , vf_active:1  },      
'{ pfvf_port:201  , pf:0 , vf:201    , vf_active:1  },      
'{ pfvf_port:202  , pf:0 , vf:202    , vf_active:1  },      
'{ pfvf_port:203  , pf:0 , vf:203    , vf_active:1  },      
'{ pfvf_port:204  , pf:0 , vf:204    , vf_active:1  },      
'{ pfvf_port:205  , pf:0 , vf:205    , vf_active:1  },      
'{ pfvf_port:206  , pf:0 , vf:206    , vf_active:1  },      
'{ pfvf_port:207  , pf:0 , vf:207    , vf_active:1  },      
'{ pfvf_port:208  , pf:0 , vf:208    , vf_active:1  },      
'{ pfvf_port:209  , pf:0 , vf:209    , vf_active:1  },      
'{ pfvf_port:210  , pf:0 , vf:210    , vf_active:1  },      
'{ pfvf_port:211  , pf:0 , vf:211    , vf_active:1  },      
'{ pfvf_port:212  , pf:0 , vf:212    , vf_active:1  },      
'{ pfvf_port:213  , pf:0 , vf:213    , vf_active:1  },      
'{ pfvf_port:214  , pf:0 , vf:214    , vf_active:1  },      
'{ pfvf_port:215  , pf:0 , vf:215    , vf_active:1  },      
'{ pfvf_port:216  , pf:0 , vf:216    , vf_active:1  },      
'{ pfvf_port:217  , pf:0 , vf:217    , vf_active:1  },      
'{ pfvf_port:218  , pf:0 , vf:218    , vf_active:1  },      
'{ pfvf_port:219  , pf:0 , vf:219    , vf_active:1  },      
'{ pfvf_port:220  , pf:0 , vf:220    , vf_active:1  },      
'{ pfvf_port:221  , pf:0 , vf:221    , vf_active:1  },      
'{ pfvf_port:222  , pf:0 , vf:222    , vf_active:1  },      
'{ pfvf_port:223  , pf:0 , vf:223    , vf_active:1  },      
'{ pfvf_port:224  , pf:0 , vf:224    , vf_active:1  },      
'{ pfvf_port:225  , pf:0 , vf:225    , vf_active:1  },      
'{ pfvf_port:226  , pf:0 , vf:226    , vf_active:1  },      
'{ pfvf_port:227  , pf:0 , vf:227    , vf_active:1  },      
'{ pfvf_port:228  , pf:0 , vf:228    , vf_active:1  },      
'{ pfvf_port:229  , pf:0 , vf:229    , vf_active:1  },      
'{ pfvf_port:230  , pf:0 , vf:230    , vf_active:1  },      
'{ pfvf_port:231  , pf:0 , vf:231    , vf_active:1  },      
'{ pfvf_port:232  , pf:0 , vf:232    , vf_active:1  },      
'{ pfvf_port:233  , pf:0 , vf:233    , vf_active:1  },      
'{ pfvf_port:234  , pf:0 , vf:234    , vf_active:1  },      
'{ pfvf_port:235  , pf:0 , vf:235    , vf_active:1  },      
'{ pfvf_port:236  , pf:0 , vf:236    , vf_active:1  },      
'{ pfvf_port:237  , pf:0 , vf:237    , vf_active:1  },      
'{ pfvf_port:238  , pf:0 , vf:238    , vf_active:1  },      
'{ pfvf_port:239  , pf:0 , vf:239    , vf_active:1  },      
'{ pfvf_port:240  , pf:0 , vf:240    , vf_active:1  },      
'{ pfvf_port:241  , pf:0 , vf:241    , vf_active:1  },      
'{ pfvf_port:242  , pf:0 , vf:242    , vf_active:1  },      
'{ pfvf_port:243  , pf:0 , vf:243    , vf_active:1  },      
'{ pfvf_port:244  , pf:0 , vf:244    , vf_active:1  },      
'{ pfvf_port:245  , pf:0 , vf:245    , vf_active:1  },      
'{ pfvf_port:246  , pf:0 , vf:246    , vf_active:1  },      
'{ pfvf_port:247  , pf:0 , vf:247    , vf_active:1  },      
'{ pfvf_port:248  , pf:0 , vf:248    , vf_active:1  },      
'{ pfvf_port:249  , pf:0 , vf:249    , vf_active:1  },      
'{ pfvf_port:250  , pf:0 , vf:250    , vf_active:1  },      
'{ pfvf_port:251  , pf:0 , vf:251    , vf_active:1  },      
'{ pfvf_port:252  , pf:0 , vf:252    , vf_active:1  },      
'{ pfvf_port:253  , pf:0 , vf:253    , vf_active:1  },      
'{ pfvf_port:254  , pf:0 , vf:254    , vf_active:1  },      
'{ pfvf_port:255  , pf:0 , vf:255    , vf_active:1  },      
'{ pfvf_port:256  , pf:0 , vf:256    , vf_active:1  },      
'{ pfvf_port:257  , pf:0 , vf:257    , vf_active:1  },      
'{ pfvf_port:258  , pf:0 , vf:258    , vf_active:1  },      
'{ pfvf_port:259  , pf:0 , vf:259    , vf_active:1  },      
'{ pfvf_port:260  , pf:0 , vf:260    , vf_active:1  },      
'{ pfvf_port:261  , pf:0 , vf:261    , vf_active:1  },      
'{ pfvf_port:262  , pf:0 , vf:262    , vf_active:1  },      
'{ pfvf_port:263  , pf:0 , vf:263    , vf_active:1  },      
'{ pfvf_port:264  , pf:0 , vf:264    , vf_active:1  },      
'{ pfvf_port:265  , pf:0 , vf:265    , vf_active:1  },      
'{ pfvf_port:266  , pf:0 , vf:266    , vf_active:1  },      
'{ pfvf_port:267  , pf:0 , vf:267    , vf_active:1  },      
'{ pfvf_port:268  , pf:0 , vf:268    , vf_active:1  },      
'{ pfvf_port:269  , pf:0 , vf:269    , vf_active:1  },      
'{ pfvf_port:270  , pf:0 , vf:270    , vf_active:1  },      
'{ pfvf_port:271  , pf:0 , vf:271    , vf_active:1  },      
'{ pfvf_port:272  , pf:0 , vf:272    , vf_active:1  },      
'{ pfvf_port:273  , pf:0 , vf:273    , vf_active:1  },      
'{ pfvf_port:274  , pf:0 , vf:274    , vf_active:1  },      
'{ pfvf_port:275  , pf:0 , vf:275    , vf_active:1  },      
'{ pfvf_port:276  , pf:0 , vf:276    , vf_active:1  },      
'{ pfvf_port:277  , pf:0 , vf:277    , vf_active:1  },      
'{ pfvf_port:278  , pf:0 , vf:278    , vf_active:1  },      
'{ pfvf_port:279  , pf:0 , vf:279    , vf_active:1  },      
'{ pfvf_port:280  , pf:0 , vf:280    , vf_active:1  },      
'{ pfvf_port:281  , pf:0 , vf:281    , vf_active:1  },      
'{ pfvf_port:282  , pf:0 , vf:282    , vf_active:1  },      
'{ pfvf_port:283  , pf:0 , vf:283    , vf_active:1  },      
'{ pfvf_port:284  , pf:0 , vf:284    , vf_active:1  },      
'{ pfvf_port:285  , pf:0 , vf:285    , vf_active:1  },      
'{ pfvf_port:286  , pf:0 , vf:286    , vf_active:1  },      
'{ pfvf_port:287  , pf:0 , vf:287    , vf_active:1  },      
'{ pfvf_port:288  , pf:0 , vf:288    , vf_active:1  },      
'{ pfvf_port:289  , pf:0 , vf:289    , vf_active:1  },      
'{ pfvf_port:290  , pf:0 , vf:290    , vf_active:1  },      
'{ pfvf_port:291  , pf:0 , vf:291    , vf_active:1  },      
'{ pfvf_port:292  , pf:0 , vf:292    , vf_active:1  },      
'{ pfvf_port:293  , pf:0 , vf:293    , vf_active:1  },      
'{ pfvf_port:294  , pf:0 , vf:294    , vf_active:1  },      
'{ pfvf_port:295  , pf:0 , vf:295    , vf_active:1  },      
'{ pfvf_port:296  , pf:0 , vf:296    , vf_active:1  },      
'{ pfvf_port:297  , pf:0 , vf:297    , vf_active:1  },      
'{ pfvf_port:298  , pf:0 , vf:298    , vf_active:1  },      
'{ pfvf_port:299  , pf:0 , vf:299    , vf_active:1  },      
'{ pfvf_port:300  , pf:0 , vf:300    , vf_active:1  },      
'{ pfvf_port:301  , pf:0 , vf:301    , vf_active:1  },      
'{ pfvf_port:302  , pf:0 , vf:302    , vf_active:1  },      
'{ pfvf_port:303  , pf:0 , vf:303    , vf_active:1  },      
'{ pfvf_port:304  , pf:0 , vf:304    , vf_active:1  },      
'{ pfvf_port:305  , pf:0 , vf:305    , vf_active:1  },      
'{ pfvf_port:306  , pf:0 , vf:306    , vf_active:1  },      
'{ pfvf_port:307  , pf:0 , vf:307    , vf_active:1  },      
'{ pfvf_port:308  , pf:0 , vf:308    , vf_active:1  },      
'{ pfvf_port:309  , pf:0 , vf:309    , vf_active:1  },      
'{ pfvf_port:310  , pf:0 , vf:310    , vf_active:1  },      
'{ pfvf_port:311  , pf:0 , vf:311    , vf_active:1  },      
'{ pfvf_port:312  , pf:0 , vf:312    , vf_active:1  },      
'{ pfvf_port:313  , pf:0 , vf:313    , vf_active:1  },      
'{ pfvf_port:314  , pf:0 , vf:314    , vf_active:1  },      
'{ pfvf_port:315  , pf:0 , vf:315    , vf_active:1  },      
'{ pfvf_port:316  , pf:0 , vf:316    , vf_active:1  },      
'{ pfvf_port:317  , pf:0 , vf:317    , vf_active:1  },      
'{ pfvf_port:318  , pf:0 , vf:318    , vf_active:1  },      
'{ pfvf_port:319  , pf:0 , vf:319    , vf_active:1  },      
'{ pfvf_port:320  , pf:0 , vf:320    , vf_active:1  },      
'{ pfvf_port:321  , pf:0 , vf:321    , vf_active:1  },      
'{ pfvf_port:322  , pf:0 , vf:322    , vf_active:1  },      
'{ pfvf_port:323  , pf:0 , vf:323    , vf_active:1  },      
'{ pfvf_port:324  , pf:0 , vf:324    , vf_active:1  },      
'{ pfvf_port:325  , pf:0 , vf:325    , vf_active:1  },      
'{ pfvf_port:326  , pf:0 , vf:326    , vf_active:1  },      
'{ pfvf_port:327  , pf:0 , vf:327    , vf_active:1  },      
'{ pfvf_port:328  , pf:0 , vf:328    , vf_active:1  },      
'{ pfvf_port:329  , pf:0 , vf:329    , vf_active:1  },      
'{ pfvf_port:330  , pf:0 , vf:330    , vf_active:1  },      
'{ pfvf_port:331  , pf:0 , vf:331    , vf_active:1  },      
'{ pfvf_port:332  , pf:0 , vf:332    , vf_active:1  },      
'{ pfvf_port:333  , pf:0 , vf:333    , vf_active:1  },      
'{ pfvf_port:334  , pf:0 , vf:334    , vf_active:1  },      
'{ pfvf_port:335  , pf:0 , vf:335    , vf_active:1  },      
'{ pfvf_port:336  , pf:0 , vf:336    , vf_active:1  },      
'{ pfvf_port:337  , pf:0 , vf:337    , vf_active:1  },      
'{ pfvf_port:338  , pf:0 , vf:338    , vf_active:1  },      
'{ pfvf_port:339  , pf:0 , vf:339    , vf_active:1  },      
'{ pfvf_port:340  , pf:0 , vf:340    , vf_active:1  },      
'{ pfvf_port:341  , pf:0 , vf:341    , vf_active:1  },      
'{ pfvf_port:342  , pf:0 , vf:342    , vf_active:1  },      
'{ pfvf_port:343  , pf:0 , vf:343    , vf_active:1  },      
'{ pfvf_port:344  , pf:0 , vf:344    , vf_active:1  },      
'{ pfvf_port:345  , pf:0 , vf:345    , vf_active:1  },      
'{ pfvf_port:346  , pf:0 , vf:346    , vf_active:1  },      
'{ pfvf_port:347  , pf:0 , vf:347    , vf_active:1  },      
'{ pfvf_port:348  , pf:0 , vf:348    , vf_active:1  },      
'{ pfvf_port:349  , pf:0 , vf:349    , vf_active:1  },      
'{ pfvf_port:350  , pf:0 , vf:350    , vf_active:1  },      
'{ pfvf_port:351  , pf:0 , vf:351    , vf_active:1  },      
'{ pfvf_port:352  , pf:0 , vf:352    , vf_active:1  },      
'{ pfvf_port:353  , pf:0 , vf:353    , vf_active:1  },      
'{ pfvf_port:354  , pf:0 , vf:354    , vf_active:1  },      
'{ pfvf_port:355  , pf:0 , vf:355    , vf_active:1  },      
'{ pfvf_port:356  , pf:0 , vf:356    , vf_active:1  },      
'{ pfvf_port:357  , pf:0 , vf:357    , vf_active:1  },      
'{ pfvf_port:358  , pf:0 , vf:358    , vf_active:1  },      
'{ pfvf_port:359  , pf:0 , vf:359    , vf_active:1  },      
'{ pfvf_port:360  , pf:0 , vf:360    , vf_active:1  },      
'{ pfvf_port:361  , pf:0 , vf:361    , vf_active:1  },      
'{ pfvf_port:362  , pf:0 , vf:362    , vf_active:1  },      
'{ pfvf_port:363  , pf:0 , vf:363    , vf_active:1  },      
'{ pfvf_port:364  , pf:0 , vf:364    , vf_active:1  },      
'{ pfvf_port:365  , pf:0 , vf:365    , vf_active:1  },      
'{ pfvf_port:366  , pf:0 , vf:366    , vf_active:1  },      
'{ pfvf_port:367  , pf:0 , vf:367    , vf_active:1  },      
'{ pfvf_port:368  , pf:0 , vf:368    , vf_active:1  },      
'{ pfvf_port:369  , pf:0 , vf:369    , vf_active:1  },      
'{ pfvf_port:370  , pf:0 , vf:370    , vf_active:1  },      
'{ pfvf_port:371  , pf:0 , vf:371    , vf_active:1  },      
'{ pfvf_port:372  , pf:0 , vf:372    , vf_active:1  },      
'{ pfvf_port:373  , pf:0 , vf:373    , vf_active:1  },      
'{ pfvf_port:374  , pf:0 , vf:374    , vf_active:1  },      
'{ pfvf_port:375  , pf:0 , vf:375    , vf_active:1  },      
'{ pfvf_port:376  , pf:0 , vf:376    , vf_active:1  },      
'{ pfvf_port:377  , pf:0 , vf:377    , vf_active:1  },      
'{ pfvf_port:378  , pf:0 , vf:378    , vf_active:1  },      
'{ pfvf_port:379  , pf:0 , vf:379    , vf_active:1  },      
'{ pfvf_port:380  , pf:0 , vf:380    , vf_active:1  },      
'{ pfvf_port:381  , pf:0 , vf:381    , vf_active:1  },      
'{ pfvf_port:382  , pf:0 , vf:382    , vf_active:1  },      
'{ pfvf_port:383  , pf:0 , vf:383    , vf_active:1  },      
'{ pfvf_port:384  , pf:0 , vf:384    , vf_active:1  },      
'{ pfvf_port:385  , pf:0 , vf:385    , vf_active:1  },      
'{ pfvf_port:386  , pf:0 , vf:386    , vf_active:1  },      
'{ pfvf_port:387  , pf:0 , vf:387    , vf_active:1  },      
'{ pfvf_port:388  , pf:0 , vf:388    , vf_active:1  },      
'{ pfvf_port:389  , pf:0 , vf:389    , vf_active:1  },      
'{ pfvf_port:390  , pf:0 , vf:390    , vf_active:1  },      
'{ pfvf_port:391  , pf:0 , vf:391    , vf_active:1  },      
'{ pfvf_port:392  , pf:0 , vf:392    , vf_active:1  },      
'{ pfvf_port:393  , pf:0 , vf:393    , vf_active:1  },      
'{ pfvf_port:394  , pf:0 , vf:394    , vf_active:1  },      
'{ pfvf_port:395  , pf:0 , vf:395    , vf_active:1  },      
'{ pfvf_port:396  , pf:0 , vf:396    , vf_active:1  },      
'{ pfvf_port:397  , pf:0 , vf:397    , vf_active:1  },      
'{ pfvf_port:398  , pf:0 , vf:398    , vf_active:1  },      
'{ pfvf_port:399  , pf:0 , vf:399    , vf_active:1  },      
'{ pfvf_port:400  , pf:0 , vf:400    , vf_active:1  },      
'{ pfvf_port:401  , pf:0 , vf:401    , vf_active:1  },      
'{ pfvf_port:402  , pf:0 , vf:402    , vf_active:1  },      
'{ pfvf_port:403  , pf:0 , vf:403    , vf_active:1  },      
'{ pfvf_port:404  , pf:0 , vf:404    , vf_active:1  },      
'{ pfvf_port:405  , pf:0 , vf:405    , vf_active:1  },      
'{ pfvf_port:406  , pf:0 , vf:406    , vf_active:1  },      
'{ pfvf_port:407  , pf:0 , vf:407    , vf_active:1  },      
'{ pfvf_port:408  , pf:0 , vf:408    , vf_active:1  },      
'{ pfvf_port:409  , pf:0 , vf:409    , vf_active:1  },      
'{ pfvf_port:410  , pf:0 , vf:410    , vf_active:1  },      
'{ pfvf_port:411  , pf:0 , vf:411    , vf_active:1  },      
'{ pfvf_port:412  , pf:0 , vf:412    , vf_active:1  },      
'{ pfvf_port:413  , pf:0 , vf:413    , vf_active:1  },      
'{ pfvf_port:414  , pf:0 , vf:414    , vf_active:1  },      
'{ pfvf_port:415  , pf:0 , vf:415    , vf_active:1  },      
'{ pfvf_port:416  , pf:0 , vf:416    , vf_active:1  },      
'{ pfvf_port:417  , pf:0 , vf:417    , vf_active:1  },      
'{ pfvf_port:418  , pf:0 , vf:418    , vf_active:1  },      
'{ pfvf_port:419  , pf:0 , vf:419    , vf_active:1  },      
'{ pfvf_port:420  , pf:0 , vf:420    , vf_active:1  },      
'{ pfvf_port:421  , pf:0 , vf:421    , vf_active:1  },      
'{ pfvf_port:422  , pf:0 , vf:422    , vf_active:1  },      
'{ pfvf_port:423  , pf:0 , vf:423    , vf_active:1  },      
'{ pfvf_port:424  , pf:0 , vf:424    , vf_active:1  },      
'{ pfvf_port:425  , pf:0 , vf:425    , vf_active:1  },      
'{ pfvf_port:426  , pf:0 , vf:426    , vf_active:1  },      
'{ pfvf_port:427  , pf:0 , vf:427    , vf_active:1  },      
'{ pfvf_port:428  , pf:0 , vf:428    , vf_active:1  },      
'{ pfvf_port:429  , pf:0 , vf:429    , vf_active:1  },      
'{ pfvf_port:430  , pf:0 , vf:430    , vf_active:1  },      
'{ pfvf_port:431  , pf:0 , vf:431    , vf_active:1  },      
'{ pfvf_port:432  , pf:0 , vf:432    , vf_active:1  },      
'{ pfvf_port:433  , pf:0 , vf:433    , vf_active:1  },      
'{ pfvf_port:434  , pf:0 , vf:434    , vf_active:1  },      
'{ pfvf_port:435  , pf:0 , vf:435    , vf_active:1  },      
'{ pfvf_port:436  , pf:0 , vf:436    , vf_active:1  },      
'{ pfvf_port:437  , pf:0 , vf:437    , vf_active:1  },      
'{ pfvf_port:438  , pf:0 , vf:438    , vf_active:1  },      
'{ pfvf_port:439  , pf:0 , vf:439    , vf_active:1  },      
'{ pfvf_port:440  , pf:0 , vf:440    , vf_active:1  },      
'{ pfvf_port:441  , pf:0 , vf:441    , vf_active:1  },      
'{ pfvf_port:442  , pf:0 , vf:442    , vf_active:1  },      
'{ pfvf_port:443  , pf:0 , vf:443    , vf_active:1  },      
'{ pfvf_port:444  , pf:0 , vf:444    , vf_active:1  },      
'{ pfvf_port:445  , pf:0 , vf:445    , vf_active:1  },      
'{ pfvf_port:446  , pf:0 , vf:446    , vf_active:1  },      
'{ pfvf_port:447  , pf:0 , vf:447    , vf_active:1  },      
'{ pfvf_port:448  , pf:0 , vf:448    , vf_active:1  },      
'{ pfvf_port:449  , pf:0 , vf:449    , vf_active:1  },
'{ pfvf_port:450  , pf:0 , vf:450    , vf_active:1  },
'{ pfvf_port:451  , pf:0 , vf:451    , vf_active:1  },
'{ pfvf_port:452  , pf:0 , vf:452    , vf_active:1  },
'{ pfvf_port:453  , pf:0 , vf:453    , vf_active:1  },
'{ pfvf_port:454  , pf:0 , vf:454    , vf_active:1  },
'{ pfvf_port:455  , pf:0 , vf:455    , vf_active:1  },
'{ pfvf_port:456  , pf:0 , vf:456    , vf_active:1  },
'{ pfvf_port:457  , pf:0 , vf:457    , vf_active:1  },
'{ pfvf_port:458  , pf:0 , vf:458    , vf_active:1  },
'{ pfvf_port:459  , pf:0 , vf:459    , vf_active:1  },
'{ pfvf_port:460  , pf:0 , vf:460    , vf_active:1  },
'{ pfvf_port:461  , pf:0 , vf:461    , vf_active:1  },
'{ pfvf_port:462  , pf:0 , vf:462    , vf_active:1  },
'{ pfvf_port:463  , pf:0 , vf:463    , vf_active:1  },
'{ pfvf_port:464  , pf:0 , vf:464    , vf_active:1  },
'{ pfvf_port:465  , pf:0 , vf:465    , vf_active:1  },
'{ pfvf_port:466  , pf:0 , vf:466    , vf_active:1  },
'{ pfvf_port:467  , pf:0 , vf:467    , vf_active:1  },
'{ pfvf_port:468  , pf:0 , vf:468    , vf_active:1  },
'{ pfvf_port:469  , pf:0 , vf:469    , vf_active:1  },
'{ pfvf_port:470  , pf:0 , vf:470    , vf_active:1  },
'{ pfvf_port:471  , pf:0 , vf:471    , vf_active:1  },
'{ pfvf_port:472  , pf:0 , vf:472    , vf_active:1  },
'{ pfvf_port:473  , pf:0 , vf:473    , vf_active:1  },
'{ pfvf_port:474  , pf:0 , vf:474    , vf_active:1  },
'{ pfvf_port:475  , pf:0 , vf:475    , vf_active:1  },
'{ pfvf_port:476  , pf:0 , vf:476    , vf_active:1  },
'{ pfvf_port:477  , pf:0 , vf:477    , vf_active:1  },
'{ pfvf_port:478  , pf:0 , vf:478    , vf_active:1  },
'{ pfvf_port:479  , pf:0 , vf:479    , vf_active:1  },
'{ pfvf_port:480  , pf:0 , vf:480    , vf_active:1  },
'{ pfvf_port:481  , pf:0 , vf:481    , vf_active:1  },
'{ pfvf_port:482  , pf:0 , vf:482    , vf_active:1  },
'{ pfvf_port:483  , pf:0 , vf:483    , vf_active:1  },
'{ pfvf_port:484  , pf:0 , vf:484    , vf_active:1  },
'{ pfvf_port:485  , pf:0 , vf:485    , vf_active:1  },
'{ pfvf_port:486  , pf:0 , vf:486    , vf_active:1  },
'{ pfvf_port:487  , pf:0 , vf:487    , vf_active:1  },
'{ pfvf_port:488  , pf:0 , vf:488    , vf_active:1  },
'{ pfvf_port:489  , pf:0 , vf:489    , vf_active:1  },
'{ pfvf_port:490  , pf:0 , vf:490    , vf_active:1  },
'{ pfvf_port:491  , pf:0 , vf:491    , vf_active:1  },
'{ pfvf_port:492  , pf:0 , vf:492    , vf_active:1  },
'{ pfvf_port:493  , pf:0 , vf:493    , vf_active:1  },
'{ pfvf_port:494  , pf:0 , vf:494    , vf_active:1  },
'{ pfvf_port:495  , pf:0 , vf:495    , vf_active:1  },
'{ pfvf_port:496  , pf:0 , vf:496    , vf_active:1  },
'{ pfvf_port:497  , pf:0 , vf:497    , vf_active:1  },
'{ pfvf_port:498  , pf:0 , vf:498    , vf_active:1  },
'{ pfvf_port:499  , pf:0 , vf:499    , vf_active:1  },
'{ pfvf_port:500  , pf:0 , vf:500    , vf_active:1  },
'{ pfvf_port:501  , pf:0 , vf:501    , vf_active:1  },
'{ pfvf_port:502  , pf:0 , vf:502    , vf_active:1  },
'{ pfvf_port:503  , pf:0 , vf:503    , vf_active:1  },
'{ pfvf_port:504  , pf:0 , vf:504    , vf_active:1  },
'{ pfvf_port:505  , pf:0 , vf:505    , vf_active:1  },
'{ pfvf_port:506  , pf:0 , vf:506    , vf_active:1  },
'{ pfvf_port:507  , pf:0 , vf:507    , vf_active:1  },
'{ pfvf_port:508  , pf:0 , vf:508    , vf_active:1  },
'{ pfvf_port:509  , pf:0 , vf:509    , vf_active:1  },
'{ pfvf_port:510  , pf:0 , vf:510    , vf_active:1  },
'{ pfvf_port:511  , pf:0 , vf:511    , vf_active:1  },
'{ pfvf_port:512  , pf:0 , vf:512    , vf_active:1  },
'{ pfvf_port:513  , pf:0 , vf:513    , vf_active:1  },
'{ pfvf_port:514  , pf:0 , vf:514    , vf_active:1  },
'{ pfvf_port:515  , pf:0 , vf:515    , vf_active:1  },
'{ pfvf_port:516  , pf:0 , vf:516    , vf_active:1  },
'{ pfvf_port:517  , pf:0 , vf:517    , vf_active:1  },
'{ pfvf_port:518  , pf:0 , vf:518    , vf_active:1  },
'{ pfvf_port:519  , pf:0 , vf:519    , vf_active:1  },
'{ pfvf_port:520  , pf:0 , vf:520    , vf_active:1  },
'{ pfvf_port:521  , pf:0 , vf:521    , vf_active:1  },
'{ pfvf_port:522  , pf:0 , vf:522    , vf_active:1  },
'{ pfvf_port:523  , pf:0 , vf:523    , vf_active:1  },
'{ pfvf_port:524  , pf:0 , vf:524    , vf_active:1  },
'{ pfvf_port:525  , pf:0 , vf:525    , vf_active:1  },
'{ pfvf_port:526  , pf:0 , vf:526    , vf_active:1  },
'{ pfvf_port:527  , pf:0 , vf:527    , vf_active:1  },
'{ pfvf_port:528  , pf:0 , vf:528    , vf_active:1  },
'{ pfvf_port:529  , pf:0 , vf:529    , vf_active:1  },
'{ pfvf_port:530  , pf:0 , vf:530    , vf_active:1  },
'{ pfvf_port:531  , pf:0 , vf:531    , vf_active:1  },
'{ pfvf_port:532  , pf:0 , vf:532    , vf_active:1  },
'{ pfvf_port:533  , pf:0 , vf:533    , vf_active:1  },
'{ pfvf_port:534  , pf:0 , vf:534    , vf_active:1  },
'{ pfvf_port:535  , pf:0 , vf:535    , vf_active:1  },
'{ pfvf_port:536  , pf:0 , vf:536    , vf_active:1  },
'{ pfvf_port:537  , pf:0 , vf:537    , vf_active:1  },
'{ pfvf_port:538  , pf:0 , vf:538    , vf_active:1  },
'{ pfvf_port:539  , pf:0 , vf:539    , vf_active:1  },
'{ pfvf_port:540  , pf:0 , vf:540    , vf_active:1  },
'{ pfvf_port:541  , pf:0 , vf:541    , vf_active:1  },
'{ pfvf_port:542  , pf:0 , vf:542    , vf_active:1  },
'{ pfvf_port:543  , pf:0 , vf:543    , vf_active:1  },
'{ pfvf_port:544  , pf:0 , vf:544    , vf_active:1  },
'{ pfvf_port:545  , pf:0 , vf:545    , vf_active:1  },
'{ pfvf_port:546  , pf:0 , vf:546    , vf_active:1  },
'{ pfvf_port:547  , pf:0 , vf:547    , vf_active:1  },
'{ pfvf_port:548  , pf:0 , vf:548    , vf_active:1  },
'{ pfvf_port:549  , pf:0 , vf:549    , vf_active:1  },
'{ pfvf_port:550  , pf:0 , vf:550    , vf_active:1  },
'{ pfvf_port:551  , pf:0 , vf:551    , vf_active:1  },
'{ pfvf_port:552  , pf:0 , vf:552    , vf_active:1  },
'{ pfvf_port:553  , pf:0 , vf:553    , vf_active:1  },
'{ pfvf_port:554  , pf:0 , vf:554    , vf_active:1  },
'{ pfvf_port:555  , pf:0 , vf:555    , vf_active:1  },
'{ pfvf_port:556  , pf:0 , vf:556    , vf_active:1  },
'{ pfvf_port:557  , pf:0 , vf:557    , vf_active:1  },
'{ pfvf_port:558  , pf:0 , vf:558    , vf_active:1  },
'{ pfvf_port:559  , pf:0 , vf:559    , vf_active:1  },
'{ pfvf_port:560  , pf:0 , vf:560    , vf_active:1  },
'{ pfvf_port:561  , pf:0 , vf:561    , vf_active:1  },
'{ pfvf_port:562  , pf:0 , vf:562    , vf_active:1  },
'{ pfvf_port:563  , pf:0 , vf:563    , vf_active:1  },
'{ pfvf_port:564  , pf:0 , vf:564    , vf_active:1  },
'{ pfvf_port:565  , pf:0 , vf:565    , vf_active:1  },
'{ pfvf_port:566  , pf:0 , vf:566    , vf_active:1  },
'{ pfvf_port:567  , pf:0 , vf:567    , vf_active:1  },
'{ pfvf_port:568  , pf:0 , vf:568    , vf_active:1  },
'{ pfvf_port:569  , pf:0 , vf:569    , vf_active:1  },
'{ pfvf_port:570  , pf:0 , vf:570    , vf_active:1  },
'{ pfvf_port:571  , pf:0 , vf:571    , vf_active:1  },
'{ pfvf_port:572  , pf:0 , vf:572    , vf_active:1  },
'{ pfvf_port:573  , pf:0 , vf:573    , vf_active:1  },
'{ pfvf_port:574  , pf:0 , vf:574    , vf_active:1  },
'{ pfvf_port:575  , pf:0 , vf:575    , vf_active:1  },
'{ pfvf_port:576  , pf:0 , vf:576    , vf_active:1  },
'{ pfvf_port:577  , pf:0 , vf:577    , vf_active:1  },
'{ pfvf_port:578  , pf:0 , vf:578    , vf_active:1  },
'{ pfvf_port:579  , pf:0 , vf:579    , vf_active:1  },
'{ pfvf_port:580  , pf:0 , vf:580    , vf_active:1  },
'{ pfvf_port:581  , pf:0 , vf:581    , vf_active:1  },
'{ pfvf_port:582  , pf:0 , vf:582    , vf_active:1  },
'{ pfvf_port:583  , pf:0 , vf:583    , vf_active:1  },
'{ pfvf_port:584  , pf:0 , vf:584    , vf_active:1  },
'{ pfvf_port:585  , pf:0 , vf:585    , vf_active:1  },
'{ pfvf_port:586  , pf:0 , vf:586    , vf_active:1  },
'{ pfvf_port:587  , pf:0 , vf:587    , vf_active:1  },
'{ pfvf_port:588  , pf:0 , vf:588    , vf_active:1  },
'{ pfvf_port:589  , pf:0 , vf:589    , vf_active:1  },
'{ pfvf_port:590  , pf:0 , vf:590    , vf_active:1  },
'{ pfvf_port:591  , pf:0 , vf:591    , vf_active:1  },
'{ pfvf_port:592  , pf:0 , vf:592    , vf_active:1  },
'{ pfvf_port:593  , pf:0 , vf:593    , vf_active:1  },
'{ pfvf_port:594  , pf:0 , vf:594    , vf_active:1  },
'{ pfvf_port:595  , pf:0 , vf:595    , vf_active:1  },
'{ pfvf_port:596  , pf:0 , vf:596    , vf_active:1  },
'{ pfvf_port:597  , pf:0 , vf:597    , vf_active:1  },
'{ pfvf_port:598  , pf:0 , vf:598    , vf_active:1  },
'{ pfvf_port:599  , pf:0 , vf:599    , vf_active:1  },
'{ pfvf_port:600  , pf:0 , vf:600    , vf_active:1  },
'{ pfvf_port:601  , pf:0 , vf:601    , vf_active:1  },
'{ pfvf_port:602  , pf:0 , vf:602    , vf_active:1  },
'{ pfvf_port:603  , pf:0 , vf:603    , vf_active:1  },
'{ pfvf_port:604  , pf:0 , vf:604    , vf_active:1  },
'{ pfvf_port:605  , pf:0 , vf:605    , vf_active:1  },
'{ pfvf_port:606  , pf:0 , vf:606    , vf_active:1  },
'{ pfvf_port:607  , pf:0 , vf:607    , vf_active:1  },
'{ pfvf_port:608  , pf:0 , vf:608    , vf_active:1  },
'{ pfvf_port:609  , pf:0 , vf:609    , vf_active:1  },
'{ pfvf_port:610  , pf:0 , vf:610    , vf_active:1  },
'{ pfvf_port:611  , pf:0 , vf:611    , vf_active:1  },
'{ pfvf_port:612  , pf:0 , vf:612    , vf_active:1  },
'{ pfvf_port:613  , pf:0 , vf:613    , vf_active:1  },
'{ pfvf_port:614  , pf:0 , vf:614    , vf_active:1  },
'{ pfvf_port:615  , pf:0 , vf:615    , vf_active:1  },
'{ pfvf_port:616  , pf:0 , vf:616    , vf_active:1  },
'{ pfvf_port:617  , pf:0 , vf:617    , vf_active:1  },
'{ pfvf_port:618  , pf:0 , vf:618    , vf_active:1  },
'{ pfvf_port:619  , pf:0 , vf:619    , vf_active:1  },
'{ pfvf_port:620  , pf:0 , vf:620    , vf_active:1  },
'{ pfvf_port:621  , pf:0 , vf:621    , vf_active:1  },
'{ pfvf_port:622  , pf:0 , vf:622    , vf_active:1  },
'{ pfvf_port:623  , pf:0 , vf:623    , vf_active:1  },
'{ pfvf_port:624  , pf:0 , vf:624    , vf_active:1  },
'{ pfvf_port:625  , pf:0 , vf:625    , vf_active:1  },
'{ pfvf_port:626  , pf:0 , vf:626    , vf_active:1  },
'{ pfvf_port:627  , pf:0 , vf:627    , vf_active:1  },
'{ pfvf_port:628  , pf:0 , vf:628    , vf_active:1  },
'{ pfvf_port:629  , pf:0 , vf:629    , vf_active:1  },
'{ pfvf_port:630  , pf:0 , vf:630    , vf_active:1  },
'{ pfvf_port:631  , pf:0 , vf:631    , vf_active:1  },
'{ pfvf_port:632  , pf:0 , vf:632    , vf_active:1  },
'{ pfvf_port:633  , pf:0 , vf:633    , vf_active:1  },
'{ pfvf_port:634  , pf:0 , vf:634    , vf_active:1  },
'{ pfvf_port:635  , pf:0 , vf:635    , vf_active:1  },
'{ pfvf_port:636  , pf:0 , vf:636    , vf_active:1  },
'{ pfvf_port:637  , pf:0 , vf:637    , vf_active:1  },
'{ pfvf_port:638  , pf:0 , vf:638    , vf_active:1  },
'{ pfvf_port:639  , pf:0 , vf:639    , vf_active:1  },
'{ pfvf_port:640  , pf:0 , vf:640    , vf_active:1  },
'{ pfvf_port:641  , pf:0 , vf:641    , vf_active:1  },
'{ pfvf_port:642  , pf:0 , vf:642    , vf_active:1  },
'{ pfvf_port:643  , pf:0 , vf:643    , vf_active:1  },
'{ pfvf_port:644  , pf:0 , vf:644    , vf_active:1  },
'{ pfvf_port:645  , pf:0 , vf:645    , vf_active:1  },
'{ pfvf_port:646  , pf:0 , vf:646    , vf_active:1  },
'{ pfvf_port:647  , pf:0 , vf:647    , vf_active:1  },
'{ pfvf_port:648  , pf:0 , vf:648    , vf_active:1  },
'{ pfvf_port:649  , pf:0 , vf:649    , vf_active:1  },
'{ pfvf_port:650  , pf:0 , vf:650    , vf_active:1  },
'{ pfvf_port:651  , pf:0 , vf:651    , vf_active:1  },
'{ pfvf_port:652  , pf:0 , vf:652    , vf_active:1  },
'{ pfvf_port:653  , pf:0 , vf:653    , vf_active:1  },
'{ pfvf_port:654  , pf:0 , vf:654    , vf_active:1  },
'{ pfvf_port:655  , pf:0 , vf:655    , vf_active:1  },
'{ pfvf_port:656  , pf:0 , vf:656    , vf_active:1  },
'{ pfvf_port:657  , pf:0 , vf:657    , vf_active:1  },
'{ pfvf_port:658  , pf:0 , vf:658    , vf_active:1  },
'{ pfvf_port:659  , pf:0 , vf:659    , vf_active:1  },
'{ pfvf_port:660  , pf:0 , vf:660    , vf_active:1  },
'{ pfvf_port:661  , pf:0 , vf:661    , vf_active:1  },
'{ pfvf_port:662  , pf:0 , vf:662    , vf_active:1  },
'{ pfvf_port:663  , pf:0 , vf:663    , vf_active:1  },
'{ pfvf_port:664  , pf:0 , vf:664    , vf_active:1  },
'{ pfvf_port:665  , pf:0 , vf:665    , vf_active:1  },
'{ pfvf_port:666  , pf:0 , vf:666    , vf_active:1  },
'{ pfvf_port:667  , pf:0 , vf:667    , vf_active:1  },
'{ pfvf_port:668  , pf:0 , vf:668    , vf_active:1  },
'{ pfvf_port:669  , pf:0 , vf:669    , vf_active:1  },
'{ pfvf_port:670  , pf:0 , vf:670    , vf_active:1  },
'{ pfvf_port:671  , pf:0 , vf:671    , vf_active:1  },
'{ pfvf_port:672  , pf:0 , vf:672    , vf_active:1  },
'{ pfvf_port:673  , pf:0 , vf:673    , vf_active:1  },
'{ pfvf_port:674  , pf:0 , vf:674    , vf_active:1  },
'{ pfvf_port:675  , pf:0 , vf:675    , vf_active:1  },
'{ pfvf_port:676  , pf:0 , vf:676    , vf_active:1  },
'{ pfvf_port:677  , pf:0 , vf:677    , vf_active:1  },
'{ pfvf_port:678  , pf:0 , vf:678    , vf_active:1  },
'{ pfvf_port:679  , pf:0 , vf:679    , vf_active:1  },
'{ pfvf_port:680  , pf:0 , vf:680    , vf_active:1  },
'{ pfvf_port:681  , pf:0 , vf:681    , vf_active:1  },
'{ pfvf_port:682  , pf:0 , vf:682    , vf_active:1  },
'{ pfvf_port:683  , pf:0 , vf:683    , vf_active:1  },
'{ pfvf_port:684  , pf:0 , vf:684    , vf_active:1  },
'{ pfvf_port:685  , pf:0 , vf:685    , vf_active:1  },
'{ pfvf_port:686  , pf:0 , vf:686    , vf_active:1  },
'{ pfvf_port:687  , pf:0 , vf:687    , vf_active:1  },
'{ pfvf_port:688  , pf:0 , vf:688    , vf_active:1  },
'{ pfvf_port:689  , pf:0 , vf:689    , vf_active:1  },
'{ pfvf_port:690  , pf:0 , vf:690    , vf_active:1  },
'{ pfvf_port:691  , pf:0 , vf:691    , vf_active:1  },
'{ pfvf_port:692  , pf:0 , vf:692    , vf_active:1  },
'{ pfvf_port:693  , pf:0 , vf:693    , vf_active:1  },
'{ pfvf_port:694  , pf:0 , vf:694    , vf_active:1  },
'{ pfvf_port:695  , pf:0 , vf:695    , vf_active:1  },
'{ pfvf_port:696  , pf:0 , vf:696    , vf_active:1  },
'{ pfvf_port:697  , pf:0 , vf:697    , vf_active:1  },
'{ pfvf_port:698  , pf:0 , vf:698    , vf_active:1  },
'{ pfvf_port:699  , pf:0 , vf:699    , vf_active:1  },
'{ pfvf_port:700  , pf:0 , vf:700    , vf_active:1  },
'{ pfvf_port:701  , pf:0 , vf:701    , vf_active:1  },
'{ pfvf_port:702  , pf:0 , vf:702    , vf_active:1  },
'{ pfvf_port:703  , pf:0 , vf:703    , vf_active:1  },
'{ pfvf_port:704  , pf:0 , vf:704    , vf_active:1  },
'{ pfvf_port:705  , pf:0 , vf:705    , vf_active:1  },
'{ pfvf_port:706  , pf:0 , vf:706    , vf_active:1  },
'{ pfvf_port:707  , pf:0 , vf:707    , vf_active:1  },
'{ pfvf_port:708  , pf:0 , vf:708    , vf_active:1  },
'{ pfvf_port:709  , pf:0 , vf:709    , vf_active:1  },
'{ pfvf_port:710  , pf:0 , vf:710    , vf_active:1  },
'{ pfvf_port:711  , pf:0 , vf:711    , vf_active:1  },
'{ pfvf_port:712  , pf:0 , vf:712    , vf_active:1  },
'{ pfvf_port:713  , pf:0 , vf:713    , vf_active:1  },
'{ pfvf_port:714  , pf:0 , vf:714    , vf_active:1  },
'{ pfvf_port:715  , pf:0 , vf:715    , vf_active:1  },
'{ pfvf_port:716  , pf:0 , vf:716    , vf_active:1  },
'{ pfvf_port:717  , pf:0 , vf:717    , vf_active:1  },
'{ pfvf_port:718  , pf:0 , vf:718    , vf_active:1  },
'{ pfvf_port:719  , pf:0 , vf:719    , vf_active:1  },
'{ pfvf_port:720  , pf:0 , vf:720    , vf_active:1  },
'{ pfvf_port:721  , pf:0 , vf:721    , vf_active:1  },
'{ pfvf_port:722  , pf:0 , vf:722    , vf_active:1  },
'{ pfvf_port:723  , pf:0 , vf:723    , vf_active:1  },
'{ pfvf_port:724  , pf:0 , vf:724    , vf_active:1  },
'{ pfvf_port:725  , pf:0 , vf:725    , vf_active:1  },
'{ pfvf_port:726  , pf:0 , vf:726    , vf_active:1  },
'{ pfvf_port:727  , pf:0 , vf:727    , vf_active:1  },
'{ pfvf_port:728  , pf:0 , vf:728    , vf_active:1  },
'{ pfvf_port:729  , pf:0 , vf:729    , vf_active:1  },
'{ pfvf_port:730  , pf:0 , vf:730    , vf_active:1  },
'{ pfvf_port:731  , pf:0 , vf:731    , vf_active:1  },
'{ pfvf_port:732  , pf:0 , vf:732    , vf_active:1  },
'{ pfvf_port:733  , pf:0 , vf:733    , vf_active:1  },
'{ pfvf_port:734  , pf:0 , vf:734    , vf_active:1  },
'{ pfvf_port:735  , pf:0 , vf:735    , vf_active:1  },
'{ pfvf_port:736  , pf:0 , vf:736    , vf_active:1  },
'{ pfvf_port:737  , pf:0 , vf:737    , vf_active:1  },
'{ pfvf_port:738  , pf:0 , vf:738    , vf_active:1  },
'{ pfvf_port:739  , pf:0 , vf:739    , vf_active:1  },
'{ pfvf_port:740  , pf:0 , vf:740    , vf_active:1  },
'{ pfvf_port:741  , pf:0 , vf:741    , vf_active:1  },
'{ pfvf_port:742  , pf:0 , vf:742    , vf_active:1  },
'{ pfvf_port:743  , pf:0 , vf:743    , vf_active:1  },
'{ pfvf_port:744  , pf:0 , vf:744    , vf_active:1  },
'{ pfvf_port:745  , pf:0 , vf:745    , vf_active:1  },
'{ pfvf_port:746  , pf:0 , vf:746    , vf_active:1  },
'{ pfvf_port:747  , pf:0 , vf:747    , vf_active:1  },
'{ pfvf_port:748  , pf:0 , vf:748    , vf_active:1  },
'{ pfvf_port:749  , pf:0 , vf:749    , vf_active:1  },
'{ pfvf_port:750  , pf:0 , vf:750    , vf_active:1  },
'{ pfvf_port:751  , pf:0 , vf:751    , vf_active:1  },
'{ pfvf_port:752  , pf:0 , vf:752    , vf_active:1  },
'{ pfvf_port:753  , pf:0 , vf:753    , vf_active:1  },
'{ pfvf_port:754  , pf:0 , vf:754    , vf_active:1  },
'{ pfvf_port:755  , pf:0 , vf:755    , vf_active:1  },
'{ pfvf_port:756  , pf:0 , vf:756    , vf_active:1  },
'{ pfvf_port:757  , pf:0 , vf:757    , vf_active:1  },
'{ pfvf_port:758  , pf:0 , vf:758    , vf_active:1  },
'{ pfvf_port:759  , pf:0 , vf:759    , vf_active:1  },
'{ pfvf_port:760  , pf:0 , vf:760    , vf_active:1  },
'{ pfvf_port:761  , pf:0 , vf:761    , vf_active:1  },
'{ pfvf_port:762  , pf:0 , vf:762    , vf_active:1  },
'{ pfvf_port:763  , pf:0 , vf:763    , vf_active:1  },
'{ pfvf_port:764  , pf:0 , vf:764    , vf_active:1  },
'{ pfvf_port:765  , pf:0 , vf:765    , vf_active:1  },
'{ pfvf_port:766  , pf:0 , vf:766    , vf_active:1  },
'{ pfvf_port:767  , pf:0 , vf:767    , vf_active:1  },
'{ pfvf_port:768  , pf:0 , vf:768    , vf_active:1  },
'{ pfvf_port:769  , pf:0 , vf:769    , vf_active:1  },
'{ pfvf_port:770  , pf:0 , vf:770    , vf_active:1  },
'{ pfvf_port:771  , pf:0 , vf:771    , vf_active:1  },
'{ pfvf_port:772  , pf:0 , vf:772    , vf_active:1  },
'{ pfvf_port:773  , pf:0 , vf:773    , vf_active:1  },
'{ pfvf_port:774  , pf:0 , vf:774    , vf_active:1  },
'{ pfvf_port:775  , pf:0 , vf:775    , vf_active:1  },
'{ pfvf_port:776  , pf:0 , vf:776    , vf_active:1  },
'{ pfvf_port:777  , pf:0 , vf:777    , vf_active:1  },
'{ pfvf_port:778  , pf:0 , vf:778    , vf_active:1  },
'{ pfvf_port:779  , pf:0 , vf:779    , vf_active:1  },
'{ pfvf_port:780  , pf:0 , vf:780    , vf_active:1  },
'{ pfvf_port:781  , pf:0 , vf:781    , vf_active:1  },
'{ pfvf_port:782  , pf:0 , vf:782    , vf_active:1  },
'{ pfvf_port:783  , pf:0 , vf:783    , vf_active:1  },
'{ pfvf_port:784  , pf:0 , vf:784    , vf_active:1  },
'{ pfvf_port:785  , pf:0 , vf:785    , vf_active:1  },
'{ pfvf_port:786  , pf:0 , vf:786    , vf_active:1  },
'{ pfvf_port:787  , pf:0 , vf:787    , vf_active:1  },
'{ pfvf_port:788  , pf:0 , vf:788    , vf_active:1  },
'{ pfvf_port:789  , pf:0 , vf:789    , vf_active:1  },
'{ pfvf_port:790  , pf:0 , vf:790    , vf_active:1  },
'{ pfvf_port:791  , pf:0 , vf:791    , vf_active:1  },
'{ pfvf_port:792  , pf:0 , vf:792    , vf_active:1  },
'{ pfvf_port:793  , pf:0 , vf:793    , vf_active:1  },
'{ pfvf_port:794  , pf:0 , vf:794    , vf_active:1  },
'{ pfvf_port:795  , pf:0 , vf:795    , vf_active:1  },
'{ pfvf_port:796  , pf:0 , vf:796    , vf_active:1  },
'{ pfvf_port:797  , pf:0 , vf:797    , vf_active:1  },
'{ pfvf_port:798  , pf:0 , vf:798    , vf_active:1  },
'{ pfvf_port:799  , pf:0 , vf:799    , vf_active:1  },
'{ pfvf_port:800  , pf:0 , vf:800    , vf_active:1  },
'{ pfvf_port:801  , pf:0 , vf:801    , vf_active:1  },
'{ pfvf_port:802  , pf:0 , vf:802    , vf_active:1  },
'{ pfvf_port:803  , pf:0 , vf:803    , vf_active:1  },
'{ pfvf_port:804  , pf:0 , vf:804    , vf_active:1  },
'{ pfvf_port:805  , pf:0 , vf:805    , vf_active:1  },
'{ pfvf_port:806  , pf:0 , vf:806    , vf_active:1  },
'{ pfvf_port:807  , pf:0 , vf:807    , vf_active:1  },
'{ pfvf_port:808  , pf:0 , vf:808    , vf_active:1  },
'{ pfvf_port:809  , pf:0 , vf:809    , vf_active:1  },
'{ pfvf_port:810  , pf:0 , vf:810    , vf_active:1  },
'{ pfvf_port:811  , pf:0 , vf:811    , vf_active:1  },
'{ pfvf_port:812  , pf:0 , vf:812    , vf_active:1  },
'{ pfvf_port:813  , pf:0 , vf:813    , vf_active:1  },
'{ pfvf_port:814  , pf:0 , vf:814    , vf_active:1  },
'{ pfvf_port:815  , pf:0 , vf:815    , vf_active:1  },
'{ pfvf_port:816  , pf:0 , vf:816    , vf_active:1  },
'{ pfvf_port:817  , pf:0 , vf:817    , vf_active:1  },
'{ pfvf_port:818  , pf:0 , vf:818    , vf_active:1  },
'{ pfvf_port:819  , pf:0 , vf:819    , vf_active:1  },
'{ pfvf_port:820  , pf:0 , vf:820    , vf_active:1  },
'{ pfvf_port:821  , pf:0 , vf:821    , vf_active:1  },
'{ pfvf_port:822  , pf:0 , vf:822    , vf_active:1  },
'{ pfvf_port:823  , pf:0 , vf:823    , vf_active:1  },
'{ pfvf_port:824  , pf:0 , vf:824    , vf_active:1  },
'{ pfvf_port:825  , pf:0 , vf:825    , vf_active:1  },
'{ pfvf_port:826  , pf:0 , vf:826    , vf_active:1  },
'{ pfvf_port:827  , pf:0 , vf:827    , vf_active:1  },
'{ pfvf_port:828  , pf:0 , vf:828    , vf_active:1  },
'{ pfvf_port:829  , pf:0 , vf:829    , vf_active:1  },
'{ pfvf_port:830  , pf:0 , vf:830    , vf_active:1  },
'{ pfvf_port:831  , pf:0 , vf:831    , vf_active:1  },
'{ pfvf_port:832  , pf:0 , vf:832    , vf_active:1  },
'{ pfvf_port:833  , pf:0 , vf:833    , vf_active:1  },
'{ pfvf_port:834  , pf:0 , vf:834    , vf_active:1  },
'{ pfvf_port:835  , pf:0 , vf:835    , vf_active:1  },
'{ pfvf_port:836  , pf:0 , vf:836    , vf_active:1  },
'{ pfvf_port:837  , pf:0 , vf:837    , vf_active:1  },
'{ pfvf_port:838  , pf:0 , vf:838    , vf_active:1  },
'{ pfvf_port:839  , pf:0 , vf:839    , vf_active:1  },
'{ pfvf_port:840  , pf:0 , vf:840    , vf_active:1  },
'{ pfvf_port:841  , pf:0 , vf:841    , vf_active:1  },
'{ pfvf_port:842  , pf:0 , vf:842    , vf_active:1  },
'{ pfvf_port:843  , pf:0 , vf:843    , vf_active:1  },
'{ pfvf_port:844  , pf:0 , vf:844    , vf_active:1  },
'{ pfvf_port:845  , pf:0 , vf:845    , vf_active:1  },
'{ pfvf_port:846  , pf:0 , vf:846    , vf_active:1  },
'{ pfvf_port:847  , pf:0 , vf:847    , vf_active:1  },
'{ pfvf_port:848  , pf:0 , vf:848    , vf_active:1  },
'{ pfvf_port:849  , pf:0 , vf:849    , vf_active:1  },
'{ pfvf_port:850  , pf:0 , vf:850    , vf_active:1  },
'{ pfvf_port:851  , pf:0 , vf:851    , vf_active:1  },
'{ pfvf_port:852  , pf:0 , vf:852    , vf_active:1  },
'{ pfvf_port:853  , pf:0 , vf:853    , vf_active:1  },
'{ pfvf_port:854  , pf:0 , vf:854    , vf_active:1  },
'{ pfvf_port:855  , pf:0 , vf:855    , vf_active:1  },
'{ pfvf_port:856  , pf:0 , vf:856    , vf_active:1  },
'{ pfvf_port:857  , pf:0 , vf:857    , vf_active:1  },
'{ pfvf_port:858  , pf:0 , vf:858    , vf_active:1  },
'{ pfvf_port:859  , pf:0 , vf:859    , vf_active:1  },
'{ pfvf_port:860  , pf:0 , vf:860    , vf_active:1  },
'{ pfvf_port:861  , pf:0 , vf:861    , vf_active:1  },
'{ pfvf_port:862  , pf:0 , vf:862    , vf_active:1  },
'{ pfvf_port:863  , pf:0 , vf:863    , vf_active:1  },
'{ pfvf_port:864  , pf:0 , vf:864    , vf_active:1  },
'{ pfvf_port:865  , pf:0 , vf:865    , vf_active:1  },
'{ pfvf_port:866  , pf:0 , vf:866    , vf_active:1  },
'{ pfvf_port:867  , pf:0 , vf:867    , vf_active:1  },
'{ pfvf_port:868  , pf:0 , vf:868    , vf_active:1  },
'{ pfvf_port:869  , pf:0 , vf:869    , vf_active:1  },
'{ pfvf_port:870  , pf:0 , vf:870    , vf_active:1  },
'{ pfvf_port:871  , pf:0 , vf:871    , vf_active:1  },
'{ pfvf_port:872  , pf:0 , vf:872    , vf_active:1  },
'{ pfvf_port:873  , pf:0 , vf:873    , vf_active:1  },
'{ pfvf_port:874  , pf:0 , vf:874    , vf_active:1  },
'{ pfvf_port:875  , pf:0 , vf:875    , vf_active:1  },
'{ pfvf_port:876  , pf:0 , vf:876    , vf_active:1  },
'{ pfvf_port:877  , pf:0 , vf:877    , vf_active:1  },
'{ pfvf_port:878  , pf:0 , vf:878    , vf_active:1  },
'{ pfvf_port:879  , pf:0 , vf:879    , vf_active:1  },
'{ pfvf_port:880  , pf:0 , vf:880    , vf_active:1  },
'{ pfvf_port:881  , pf:0 , vf:881    , vf_active:1  },
'{ pfvf_port:882  , pf:0 , vf:882    , vf_active:1  },
'{ pfvf_port:883  , pf:0 , vf:883    , vf_active:1  },
'{ pfvf_port:884  , pf:0 , vf:884    , vf_active:1  },
'{ pfvf_port:885  , pf:0 , vf:885    , vf_active:1  },
'{ pfvf_port:886  , pf:0 , vf:886    , vf_active:1  },
'{ pfvf_port:887  , pf:0 , vf:887    , vf_active:1  },
'{ pfvf_port:888  , pf:0 , vf:888    , vf_active:1  },
'{ pfvf_port:889  , pf:0 , vf:889    , vf_active:1  },
'{ pfvf_port:890  , pf:0 , vf:890    , vf_active:1  },
'{ pfvf_port:891  , pf:0 , vf:891    , vf_active:1  },
'{ pfvf_port:892  , pf:0 , vf:892    , vf_active:1  },
'{ pfvf_port:893  , pf:0 , vf:893    , vf_active:1  },
'{ pfvf_port:894  , pf:0 , vf:894    , vf_active:1  },
'{ pfvf_port:895  , pf:0 , vf:895    , vf_active:1  },
'{ pfvf_port:896  , pf:0 , vf:896    , vf_active:1  },
'{ pfvf_port:897  , pf:0 , vf:897    , vf_active:1  },
'{ pfvf_port:898  , pf:0 , vf:898    , vf_active:1  },
'{ pfvf_port:899  , pf:0 , vf:899    , vf_active:1  },
'{ pfvf_port:900  , pf:0 , vf:900    , vf_active:1  },
'{ pfvf_port:901  , pf:0 , vf:901    , vf_active:1  },
'{ pfvf_port:902  , pf:0 , vf:902    , vf_active:1  },
'{ pfvf_port:903  , pf:0 , vf:903    , vf_active:1  },
'{ pfvf_port:904  , pf:0 , vf:904    , vf_active:1  },
'{ pfvf_port:905  , pf:0 , vf:905    , vf_active:1  },
'{ pfvf_port:906  , pf:0 , vf:906    , vf_active:1  },
'{ pfvf_port:907  , pf:0 , vf:907    , vf_active:1  },
'{ pfvf_port:908  , pf:0 , vf:908    , vf_active:1  },
'{ pfvf_port:909  , pf:0 , vf:909    , vf_active:1  },
'{ pfvf_port:910  , pf:0 , vf:910    , vf_active:1  },
'{ pfvf_port:911  , pf:0 , vf:911    , vf_active:1  },
'{ pfvf_port:912  , pf:0 , vf:912    , vf_active:1  },
'{ pfvf_port:913  , pf:0 , vf:913    , vf_active:1  },
'{ pfvf_port:914  , pf:0 , vf:914    , vf_active:1  },
'{ pfvf_port:915  , pf:0 , vf:915    , vf_active:1  },
'{ pfvf_port:916  , pf:0 , vf:916    , vf_active:1  },
'{ pfvf_port:917  , pf:0 , vf:917    , vf_active:1  },
'{ pfvf_port:918  , pf:0 , vf:918    , vf_active:1  },
'{ pfvf_port:919  , pf:0 , vf:919    , vf_active:1  },
'{ pfvf_port:920  , pf:0 , vf:920    , vf_active:1  },
'{ pfvf_port:921  , pf:0 , vf:921    , vf_active:1  },
'{ pfvf_port:922  , pf:0 , vf:922    , vf_active:1  },
'{ pfvf_port:923  , pf:0 , vf:923    , vf_active:1  },
'{ pfvf_port:924  , pf:0 , vf:924    , vf_active:1  },
'{ pfvf_port:925  , pf:0 , vf:925    , vf_active:1  },
'{ pfvf_port:926  , pf:0 , vf:926    , vf_active:1  },
'{ pfvf_port:927  , pf:0 , vf:927    , vf_active:1  },
'{ pfvf_port:928  , pf:0 , vf:928    , vf_active:1  },
'{ pfvf_port:929  , pf:0 , vf:929    , vf_active:1  },
'{ pfvf_port:930  , pf:0 , vf:930    , vf_active:1  },
'{ pfvf_port:931  , pf:0 , vf:931    , vf_active:1  },
'{ pfvf_port:932  , pf:0 , vf:932    , vf_active:1  },
'{ pfvf_port:933  , pf:0 , vf:933    , vf_active:1  },
'{ pfvf_port:934  , pf:0 , vf:934    , vf_active:1  },
'{ pfvf_port:935  , pf:0 , vf:935    , vf_active:1  },
'{ pfvf_port:936  , pf:0 , vf:936    , vf_active:1  },
'{ pfvf_port:937  , pf:0 , vf:937    , vf_active:1  },
'{ pfvf_port:938  , pf:0 , vf:938    , vf_active:1  },
'{ pfvf_port:939  , pf:0 , vf:939    , vf_active:1  },
'{ pfvf_port:940  , pf:0 , vf:940    , vf_active:1  },
'{ pfvf_port:941  , pf:0 , vf:941    , vf_active:1  },
'{ pfvf_port:942  , pf:0 , vf:942    , vf_active:1  },
'{ pfvf_port:943  , pf:0 , vf:943    , vf_active:1  },
'{ pfvf_port:944  , pf:0 , vf:944    , vf_active:1  },
'{ pfvf_port:945  , pf:0 , vf:945    , vf_active:1  },
'{ pfvf_port:946  , pf:0 , vf:946    , vf_active:1  },
'{ pfvf_port:947  , pf:0 , vf:947    , vf_active:1  },
'{ pfvf_port:948  , pf:0 , vf:948    , vf_active:1  },
'{ pfvf_port:949  , pf:0 , vf:949    , vf_active:1  },
'{ pfvf_port:950  , pf:0 , vf:950    , vf_active:1  },
'{ pfvf_port:951  , pf:0 , vf:951    , vf_active:1  },
'{ pfvf_port:952  , pf:0 , vf:952    , vf_active:1  },
'{ pfvf_port:953  , pf:0 , vf:953    , vf_active:1  },
'{ pfvf_port:954  , pf:0 , vf:954    , vf_active:1  },
'{ pfvf_port:955  , pf:0 , vf:955    , vf_active:1  },
'{ pfvf_port:956  , pf:0 , vf:956    , vf_active:1  },
'{ pfvf_port:957  , pf:0 , vf:957    , vf_active:1  },
'{ pfvf_port:958  , pf:0 , vf:958    , vf_active:1  },
'{ pfvf_port:959  , pf:0 , vf:959    , vf_active:1  },
'{ pfvf_port:960  , pf:0 , vf:960    , vf_active:1  },
'{ pfvf_port:961  , pf:0 , vf:961    , vf_active:1  },
'{ pfvf_port:962  , pf:0 , vf:962    , vf_active:1  },
'{ pfvf_port:963  , pf:0 , vf:963    , vf_active:1  },
'{ pfvf_port:964  , pf:0 , vf:964    , vf_active:1  },
'{ pfvf_port:965  , pf:0 , vf:965    , vf_active:1  },
'{ pfvf_port:966  , pf:0 , vf:966    , vf_active:1  },
'{ pfvf_port:967  , pf:0 , vf:967    , vf_active:1  },
'{ pfvf_port:968  , pf:0 , vf:968    , vf_active:1  },
'{ pfvf_port:969  , pf:0 , vf:969    , vf_active:1  },
'{ pfvf_port:970  , pf:0 , vf:970    , vf_active:1  },
'{ pfvf_port:971  , pf:0 , vf:971    , vf_active:1  },
'{ pfvf_port:972  , pf:0 , vf:972    , vf_active:1  },
'{ pfvf_port:973  , pf:0 , vf:973    , vf_active:1  },
'{ pfvf_port:974  , pf:0 , vf:974    , vf_active:1  },
'{ pfvf_port:975  , pf:0 , vf:975    , vf_active:1  },
'{ pfvf_port:976  , pf:0 , vf:976    , vf_active:1  },
'{ pfvf_port:977  , pf:0 , vf:977    , vf_active:1  },
'{ pfvf_port:978  , pf:0 , vf:978    , vf_active:1  },
'{ pfvf_port:979  , pf:0 , vf:979    , vf_active:1  },
'{ pfvf_port:980  , pf:0 , vf:980    , vf_active:1  },
'{ pfvf_port:981  , pf:0 , vf:981    , vf_active:1  },
'{ pfvf_port:982  , pf:0 , vf:982    , vf_active:1  },
'{ pfvf_port:983  , pf:0 , vf:983    , vf_active:1  },
'{ pfvf_port:984  , pf:0 , vf:984    , vf_active:1  },
'{ pfvf_port:985  , pf:0 , vf:985    , vf_active:1  },
'{ pfvf_port:986  , pf:0 , vf:986    , vf_active:1  },
'{ pfvf_port:987  , pf:0 , vf:987    , vf_active:1  },
'{ pfvf_port:988  , pf:0 , vf:988    , vf_active:1  },
'{ pfvf_port:989  , pf:0 , vf:989    , vf_active:1  },
'{ pfvf_port:990  , pf:0 , vf:990    , vf_active:1  },
'{ pfvf_port:991  , pf:0 , vf:991    , vf_active:1  },
'{ pfvf_port:992  , pf:0 , vf:992    , vf_active:1  },
'{ pfvf_port:993  , pf:0 , vf:993    , vf_active:1  },
'{ pfvf_port:994  , pf:0 , vf:994    , vf_active:1  },
'{ pfvf_port:995  , pf:0 , vf:995    , vf_active:1  },
'{ pfvf_port:996  , pf:0 , vf:996    , vf_active:1  },
'{ pfvf_port:997  , pf:0 , vf:997    , vf_active:1  },
'{ pfvf_port:998  , pf:0 , vf:998    , vf_active:1  },
'{ pfvf_port:999  , pf:0 , vf:999    , vf_active:1  },
'{ pfvf_port:1000  , pf:0 , vf:1000    , vf_active:1  },
'{ pfvf_port:1001  , pf:0 , vf:1001    , vf_active:1  },
'{ pfvf_port:1002  , pf:0 , vf:1002    , vf_active:1  },
'{ pfvf_port:1003  , pf:0 , vf:1003    , vf_active:1  },
'{ pfvf_port:1004  , pf:0 , vf:1004    , vf_active:1  },
'{ pfvf_port:1005  , pf:0 , vf:1005    , vf_active:1  },
'{ pfvf_port:1006  , pf:0 , vf:1006    , vf_active:1  },
'{ pfvf_port:1007  , pf:0 , vf:1007    , vf_active:1  },
'{ pfvf_port:1008  , pf:0 , vf:1008    , vf_active:1  },
'{ pfvf_port:1009  , pf:0 , vf:1009    , vf_active:1  },
'{ pfvf_port:1010  , pf:0 , vf:1010    , vf_active:1  },
'{ pfvf_port:1011  , pf:0 , vf:1011    , vf_active:1  },
'{ pfvf_port:1012  , pf:0 , vf:1012    , vf_active:1  },
'{ pfvf_port:1013  , pf:0 , vf:1013    , vf_active:1  },
'{ pfvf_port:1014  , pf:0 , vf:1014    , vf_active:1  },
'{ pfvf_port:1015  , pf:0 , vf:1015    , vf_active:1  },
'{ pfvf_port:1016  , pf:0 , vf:1016    , vf_active:1  },
'{ pfvf_port:1017  , pf:0 , vf:1017    , vf_active:1  },
'{ pfvf_port:1018  , pf:0 , vf:1018    , vf_active:1  },
'{ pfvf_port:1019  , pf:0 , vf:1019    , vf_active:1  },
'{ pfvf_port:1020  , pf:0 , vf:1020    , vf_active:1  },
'{ pfvf_port:1021  , pf:0 , vf:1021    , vf_active:1  },
'{ pfvf_port:1022  , pf:0 , vf:1022    , vf_active:1  },
'{ pfvf_port:1023  , pf:0 , vf:1023    , vf_active:1  },
'{ pfvf_port:1024  , pf:0 , vf:1024    , vf_active:1  },
'{ pfvf_port:1025  , pf:0 , vf:1025    , vf_active:1  },
'{ pfvf_port:1026  , pf:0 , vf:1026    , vf_active:1  },
'{ pfvf_port:1027  , pf:0 , vf:1027    , vf_active:1  },
'{ pfvf_port:1028  , pf:0 , vf:1028    , vf_active:1  },
'{ pfvf_port:1029  , pf:0 , vf:1029    , vf_active:1  },
'{ pfvf_port:1030  , pf:0 , vf:1030    , vf_active:1  },
'{ pfvf_port:1031  , pf:0 , vf:1031    , vf_active:1  },
'{ pfvf_port:1032  , pf:0 , vf:1032    , vf_active:1  },
'{ pfvf_port:1033  , pf:0 , vf:1033    , vf_active:1  },
'{ pfvf_port:1034  , pf:0 , vf:1034    , vf_active:1  },
'{ pfvf_port:1035  , pf:0 , vf:1035    , vf_active:1  },
'{ pfvf_port:1036  , pf:0 , vf:1036    , vf_active:1  },
'{ pfvf_port:1037  , pf:0 , vf:1037    , vf_active:1  },
'{ pfvf_port:1038  , pf:0 , vf:1038    , vf_active:1  },
'{ pfvf_port:1039  , pf:0 , vf:1039    , vf_active:1  },
'{ pfvf_port:1040  , pf:0 , vf:1040    , vf_active:1  },
'{ pfvf_port:1041  , pf:0 , vf:1041    , vf_active:1  },
'{ pfvf_port:1042  , pf:0 , vf:1042    , vf_active:1  },
'{ pfvf_port:1043  , pf:0 , vf:1043    , vf_active:1  },
'{ pfvf_port:1044  , pf:0 , vf:1044    , vf_active:1  },
'{ pfvf_port:1045  , pf:0 , vf:1045    , vf_active:1  },
'{ pfvf_port:1046  , pf:0 , vf:1046    , vf_active:1  },
'{ pfvf_port:1047  , pf:0 , vf:1047    , vf_active:1  },
'{ pfvf_port:1048  , pf:0 , vf:1048    , vf_active:1  },
'{ pfvf_port:1049  , pf:0 , vf:1049    , vf_active:1  },
'{ pfvf_port:1050  , pf:0 , vf:1050    , vf_active:1  },
'{ pfvf_port:1051  , pf:0 , vf:1051    , vf_active:1  },
'{ pfvf_port:1052  , pf:0 , vf:1052    , vf_active:1  },
'{ pfvf_port:1053  , pf:0 , vf:1053    , vf_active:1  },
'{ pfvf_port:1054  , pf:0 , vf:1054    , vf_active:1  },
'{ pfvf_port:1055  , pf:0 , vf:1055    , vf_active:1  },
'{ pfvf_port:1056  , pf:0 , vf:1056    , vf_active:1  },
'{ pfvf_port:1057  , pf:0 , vf:1057    , vf_active:1  },
'{ pfvf_port:1058  , pf:0 , vf:1058    , vf_active:1  },
'{ pfvf_port:1059  , pf:0 , vf:1059    , vf_active:1  },
'{ pfvf_port:1060  , pf:0 , vf:1060    , vf_active:1  },
'{ pfvf_port:1061  , pf:0 , vf:1061    , vf_active:1  },
'{ pfvf_port:1062  , pf:0 , vf:1062    , vf_active:1  },
'{ pfvf_port:1063  , pf:0 , vf:1063    , vf_active:1  },
'{ pfvf_port:1064  , pf:0 , vf:1064    , vf_active:1  },
'{ pfvf_port:1065  , pf:0 , vf:1065    , vf_active:1  },
'{ pfvf_port:1066  , pf:0 , vf:1066    , vf_active:1  },
'{ pfvf_port:1067  , pf:0 , vf:1067    , vf_active:1  },
'{ pfvf_port:1068  , pf:0 , vf:1068    , vf_active:1  },
'{ pfvf_port:1069  , pf:0 , vf:1069    , vf_active:1  },
'{ pfvf_port:1070  , pf:0 , vf:1070    , vf_active:1  },
'{ pfvf_port:1071  , pf:0 , vf:1071    , vf_active:1  },
'{ pfvf_port:1072  , pf:0 , vf:1072    , vf_active:1  },
'{ pfvf_port:1073  , pf:0 , vf:1073    , vf_active:1  },
'{ pfvf_port:1074  , pf:0 , vf:1074    , vf_active:1  },
'{ pfvf_port:1075  , pf:0 , vf:1075    , vf_active:1  },
'{ pfvf_port:1076  , pf:0 , vf:1076    , vf_active:1  },
'{ pfvf_port:1077  , pf:0 , vf:1077    , vf_active:1  },
'{ pfvf_port:1078  , pf:0 , vf:1078    , vf_active:1  },
'{ pfvf_port:1079  , pf:0 , vf:1079    , vf_active:1  },
'{ pfvf_port:1080  , pf:0 , vf:1080    , vf_active:1  },
'{ pfvf_port:1081  , pf:0 , vf:1081    , vf_active:1  },
'{ pfvf_port:1082  , pf:0 , vf:1082    , vf_active:1  },
'{ pfvf_port:1083  , pf:0 , vf:1083    , vf_active:1  },
'{ pfvf_port:1084  , pf:0 , vf:1084    , vf_active:1  },
'{ pfvf_port:1085  , pf:0 , vf:1085    , vf_active:1  },
'{ pfvf_port:1086  , pf:0 , vf:1086    , vf_active:1  },
'{ pfvf_port:1087  , pf:0 , vf:1087    , vf_active:1  },
'{ pfvf_port:1088  , pf:0 , vf:1088    , vf_active:1  },
'{ pfvf_port:1089  , pf:0 , vf:1089    , vf_active:1  },
'{ pfvf_port:1090  , pf:0 , vf:1090    , vf_active:1  },
'{ pfvf_port:1091  , pf:0 , vf:1091    , vf_active:1  },
'{ pfvf_port:1092  , pf:0 , vf:1092    , vf_active:1  },
'{ pfvf_port:1093  , pf:0 , vf:1093    , vf_active:1  },
'{ pfvf_port:1094  , pf:0 , vf:1094    , vf_active:1  },
'{ pfvf_port:1095  , pf:0 , vf:1095    , vf_active:1  },
'{ pfvf_port:1096  , pf:0 , vf:1096    , vf_active:1  },
'{ pfvf_port:1097  , pf:0 , vf:1097    , vf_active:1  },
'{ pfvf_port:1098  , pf:0 , vf:1098    , vf_active:1  },
'{ pfvf_port:1099  , pf:0 , vf:1099    , vf_active:1  },
'{ pfvf_port:1100  , pf:0 , vf:1100    , vf_active:1  },
'{ pfvf_port:1101  , pf:0 , vf:1101    , vf_active:1  },
'{ pfvf_port:1102  , pf:0 , vf:1102    , vf_active:1  },
'{ pfvf_port:1103  , pf:0 , vf:1103    , vf_active:1  },
'{ pfvf_port:1104  , pf:0 , vf:1104    , vf_active:1  },
'{ pfvf_port:1105  , pf:0 , vf:1105    , vf_active:1  },
'{ pfvf_port:1106  , pf:0 , vf:1106    , vf_active:1  },
'{ pfvf_port:1107  , pf:0 , vf:1107    , vf_active:1  },
'{ pfvf_port:1108  , pf:0 , vf:1108    , vf_active:1  },
'{ pfvf_port:1109  , pf:0 , vf:1109    , vf_active:1  },
'{ pfvf_port:1110  , pf:0 , vf:1110    , vf_active:1  },
'{ pfvf_port:1111  , pf:0 , vf:1111    , vf_active:1  },
'{ pfvf_port:1112  , pf:0 , vf:1112    , vf_active:1  },
'{ pfvf_port:1113  , pf:0 , vf:1113    , vf_active:1  },
'{ pfvf_port:1114  , pf:0 , vf:1114    , vf_active:1  },
'{ pfvf_port:1115  , pf:0 , vf:1115    , vf_active:1  },
'{ pfvf_port:1116  , pf:0 , vf:1116    , vf_active:1  },
'{ pfvf_port:1117  , pf:0 , vf:1117    , vf_active:1  },
'{ pfvf_port:1118  , pf:0 , vf:1118    , vf_active:1  },
'{ pfvf_port:1119  , pf:0 , vf:1119    , vf_active:1  },
'{ pfvf_port:1120  , pf:0 , vf:1120    , vf_active:1  },
'{ pfvf_port:1121  , pf:0 , vf:1121    , vf_active:1  },
'{ pfvf_port:1122  , pf:0 , vf:1122    , vf_active:1  },
'{ pfvf_port:1123  , pf:0 , vf:1123    , vf_active:1  },
'{ pfvf_port:1124  , pf:0 , vf:1124    , vf_active:1  },
'{ pfvf_port:1125  , pf:0 , vf:1125    , vf_active:1  },
'{ pfvf_port:1126  , pf:0 , vf:1126    , vf_active:1  },
'{ pfvf_port:1127  , pf:0 , vf:1127    , vf_active:1  },
'{ pfvf_port:1128  , pf:0 , vf:1128    , vf_active:1  },
'{ pfvf_port:1129  , pf:0 , vf:1129    , vf_active:1  },
'{ pfvf_port:1130  , pf:0 , vf:1130    , vf_active:1  },
'{ pfvf_port:1131  , pf:0 , vf:1131    , vf_active:1  },
'{ pfvf_port:1132  , pf:0 , vf:1132    , vf_active:1  },
'{ pfvf_port:1133  , pf:0 , vf:1133    , vf_active:1  },
'{ pfvf_port:1134  , pf:0 , vf:1134    , vf_active:1  },
'{ pfvf_port:1135  , pf:0 , vf:1135    , vf_active:1  },
'{ pfvf_port:1136  , pf:0 , vf:1136    , vf_active:1  },
'{ pfvf_port:1137  , pf:0 , vf:1137    , vf_active:1  },
'{ pfvf_port:1138  , pf:0 , vf:1138    , vf_active:1  },
'{ pfvf_port:1139  , pf:0 , vf:1139    , vf_active:1  },
'{ pfvf_port:1140  , pf:0 , vf:1140    , vf_active:1  },
'{ pfvf_port:1141  , pf:0 , vf:1141    , vf_active:1  },
'{ pfvf_port:1142  , pf:0 , vf:1142    , vf_active:1  },
'{ pfvf_port:1143  , pf:0 , vf:1143    , vf_active:1  },
'{ pfvf_port:1144  , pf:0 , vf:1144    , vf_active:1  },
'{ pfvf_port:1145  , pf:0 , vf:1145    , vf_active:1  },
'{ pfvf_port:1146  , pf:0 , vf:1146    , vf_active:1  },
'{ pfvf_port:1147  , pf:0 , vf:1147    , vf_active:1  },
'{ pfvf_port:1148  , pf:0 , vf:1148    , vf_active:1  },
'{ pfvf_port:1149  , pf:0 , vf:1149    , vf_active:1  },
'{ pfvf_port:1150  , pf:0 , vf:1150    , vf_active:1  },
'{ pfvf_port:1151  , pf:0 , vf:1151    , vf_active:1  },
'{ pfvf_port:1152  , pf:0 , vf:1152    , vf_active:1  },
'{ pfvf_port:1153  , pf:0 , vf:1153    , vf_active:1  },
'{ pfvf_port:1154  , pf:0 , vf:1154    , vf_active:1  },
'{ pfvf_port:1155  , pf:0 , vf:1155    , vf_active:1  },
'{ pfvf_port:1156  , pf:0 , vf:1156    , vf_active:1  },
'{ pfvf_port:1157  , pf:0 , vf:1157    , vf_active:1  },
'{ pfvf_port:1158  , pf:0 , vf:1158    , vf_active:1  },
'{ pfvf_port:1159  , pf:0 , vf:1159    , vf_active:1  },
'{ pfvf_port:1160  , pf:0 , vf:1160    , vf_active:1  },
'{ pfvf_port:1161  , pf:0 , vf:1161    , vf_active:1  },
'{ pfvf_port:1162  , pf:0 , vf:1162    , vf_active:1  },
'{ pfvf_port:1163  , pf:0 , vf:1163    , vf_active:1  },
'{ pfvf_port:1164  , pf:0 , vf:1164    , vf_active:1  },
'{ pfvf_port:1165  , pf:0 , vf:1165    , vf_active:1  },
'{ pfvf_port:1166  , pf:0 , vf:1166    , vf_active:1  },
'{ pfvf_port:1167  , pf:0 , vf:1167    , vf_active:1  },
'{ pfvf_port:1168  , pf:0 , vf:1168    , vf_active:1  },
'{ pfvf_port:1169  , pf:0 , vf:1169    , vf_active:1  },
'{ pfvf_port:1170  , pf:0 , vf:1170    , vf_active:1  },
'{ pfvf_port:1171  , pf:0 , vf:1171    , vf_active:1  },
'{ pfvf_port:1172  , pf:0 , vf:1172    , vf_active:1  },
'{ pfvf_port:1173  , pf:0 , vf:1173    , vf_active:1  },
'{ pfvf_port:1174  , pf:0 , vf:1174    , vf_active:1  },
'{ pfvf_port:1175  , pf:0 , vf:1175    , vf_active:1  },
'{ pfvf_port:1176  , pf:0 , vf:1176    , vf_active:1  },
'{ pfvf_port:1177  , pf:0 , vf:1177    , vf_active:1  },
'{ pfvf_port:1178  , pf:0 , vf:1178    , vf_active:1  },
'{ pfvf_port:1179  , pf:0 , vf:1179    , vf_active:1  },
'{ pfvf_port:1180  , pf:0 , vf:1180    , vf_active:1  },
'{ pfvf_port:1181  , pf:0 , vf:1181    , vf_active:1  },
'{ pfvf_port:1182  , pf:0 , vf:1182    , vf_active:1  },
'{ pfvf_port:1183  , pf:0 , vf:1183    , vf_active:1  },
'{ pfvf_port:1184  , pf:0 , vf:1184    , vf_active:1  },
'{ pfvf_port:1185  , pf:0 , vf:1185    , vf_active:1  },
'{ pfvf_port:1186  , pf:0 , vf:1186    , vf_active:1  },
'{ pfvf_port:1187  , pf:0 , vf:1187    , vf_active:1  },
'{ pfvf_port:1188  , pf:0 , vf:1188    , vf_active:1  },
'{ pfvf_port:1189  , pf:0 , vf:1189    , vf_active:1  },
'{ pfvf_port:1190  , pf:0 , vf:1190    , vf_active:1  },
'{ pfvf_port:1191  , pf:0 , vf:1191    , vf_active:1  },
'{ pfvf_port:1192  , pf:0 , vf:1192    , vf_active:1  },
'{ pfvf_port:1193  , pf:0 , vf:1193    , vf_active:1  },
'{ pfvf_port:1194  , pf:0 , vf:1194    , vf_active:1  },
'{ pfvf_port:1195  , pf:0 , vf:1195    , vf_active:1  },
'{ pfvf_port:1196  , pf:0 , vf:1196    , vf_active:1  },
'{ pfvf_port:1197  , pf:0 , vf:1197    , vf_active:1  },
'{ pfvf_port:1198  , pf:0 , vf:1198    , vf_active:1  },
'{ pfvf_port:1199  , pf:0 , vf:1199    , vf_active:1  },
'{ pfvf_port:1200  , pf:0 , vf:1200    , vf_active:1  },
'{ pfvf_port:1201  , pf:0 , vf:1201    , vf_active:1  },
'{ pfvf_port:1202  , pf:0 , vf:1202    , vf_active:1  },
'{ pfvf_port:1203  , pf:0 , vf:1203    , vf_active:1  },
'{ pfvf_port:1204  , pf:0 , vf:1204    , vf_active:1  },
'{ pfvf_port:1205  , pf:0 , vf:1205    , vf_active:1  },
'{ pfvf_port:1206  , pf:0 , vf:1206    , vf_active:1  },
'{ pfvf_port:1207  , pf:0 , vf:1207    , vf_active:1  },
'{ pfvf_port:1208  , pf:0 , vf:1208    , vf_active:1  },
'{ pfvf_port:1209  , pf:0 , vf:1209    , vf_active:1  },
'{ pfvf_port:1210  , pf:0 , vf:1210    , vf_active:1  },
'{ pfvf_port:1211  , pf:0 , vf:1211    , vf_active:1  },
'{ pfvf_port:1212  , pf:0 , vf:1212    , vf_active:1  },
'{ pfvf_port:1213  , pf:0 , vf:1213    , vf_active:1  },
'{ pfvf_port:1214  , pf:0 , vf:1214    , vf_active:1  },
'{ pfvf_port:1215  , pf:0 , vf:1215    , vf_active:1  },
'{ pfvf_port:1216  , pf:0 , vf:1216    , vf_active:1  },
'{ pfvf_port:1217  , pf:0 , vf:1217    , vf_active:1  },
'{ pfvf_port:1218  , pf:0 , vf:1218    , vf_active:1  },
'{ pfvf_port:1219  , pf:0 , vf:1219    , vf_active:1  },
'{ pfvf_port:1220  , pf:0 , vf:1220    , vf_active:1  },
'{ pfvf_port:1221  , pf:0 , vf:1221    , vf_active:1  },
'{ pfvf_port:1222  , pf:0 , vf:1222    , vf_active:1  },
'{ pfvf_port:1223  , pf:0 , vf:1223    , vf_active:1  },
'{ pfvf_port:1224  , pf:0 , vf:1224    , vf_active:1  },
'{ pfvf_port:1225  , pf:0 , vf:1225    , vf_active:1  },
'{ pfvf_port:1226  , pf:0 , vf:1226    , vf_active:1  },
'{ pfvf_port:1227  , pf:0 , vf:1227    , vf_active:1  },
'{ pfvf_port:1228  , pf:0 , vf:1228    , vf_active:1  },
'{ pfvf_port:1229  , pf:0 , vf:1229    , vf_active:1  },
'{ pfvf_port:1230  , pf:0 , vf:1230    , vf_active:1  },
'{ pfvf_port:1231  , pf:0 , vf:1231    , vf_active:1  },
'{ pfvf_port:1232  , pf:0 , vf:1232    , vf_active:1  },
'{ pfvf_port:1233  , pf:0 , vf:1233    , vf_active:1  },
'{ pfvf_port:1234  , pf:0 , vf:1234    , vf_active:1  },
'{ pfvf_port:1235  , pf:0 , vf:1235    , vf_active:1  },
'{ pfvf_port:1236  , pf:0 , vf:1236    , vf_active:1  },
'{ pfvf_port:1237  , pf:0 , vf:1237    , vf_active:1  },
'{ pfvf_port:1238  , pf:0 , vf:1238    , vf_active:1  },
'{ pfvf_port:1239  , pf:0 , vf:1239    , vf_active:1  },
'{ pfvf_port:1240  , pf:0 , vf:1240    , vf_active:1  },
'{ pfvf_port:1241  , pf:0 , vf:1241    , vf_active:1  },
'{ pfvf_port:1242  , pf:0 , vf:1242    , vf_active:1  },
'{ pfvf_port:1243  , pf:0 , vf:1243    , vf_active:1  },
'{ pfvf_port:1244  , pf:0 , vf:1244    , vf_active:1  },
'{ pfvf_port:1245  , pf:0 , vf:1245    , vf_active:1  },
'{ pfvf_port:1246  , pf:0 , vf:1246    , vf_active:1  },
'{ pfvf_port:1247  , pf:0 , vf:1247    , vf_active:1  },
'{ pfvf_port:1248  , pf:0 , vf:1248    , vf_active:1  },
'{ pfvf_port:1249  , pf:0 , vf:1249    , vf_active:1  },
'{ pfvf_port:1250  , pf:0 , vf:1250    , vf_active:1  },
'{ pfvf_port:1251  , pf:0 , vf:1251    , vf_active:1  },
'{ pfvf_port:1252  , pf:0 , vf:1252    , vf_active:1  },
'{ pfvf_port:1253  , pf:0 , vf:1253    , vf_active:1  },
'{ pfvf_port:1254  , pf:0 , vf:1254    , vf_active:1  },
'{ pfvf_port:1255  , pf:0 , vf:1255    , vf_active:1  },
'{ pfvf_port:1256  , pf:0 , vf:1256    , vf_active:1  },
'{ pfvf_port:1257  , pf:0 , vf:1257    , vf_active:1  },
'{ pfvf_port:1258  , pf:0 , vf:1258    , vf_active:1  },
'{ pfvf_port:1259  , pf:0 , vf:1259    , vf_active:1  },
'{ pfvf_port:1260  , pf:0 , vf:1260    , vf_active:1  },
'{ pfvf_port:1261  , pf:0 , vf:1261    , vf_active:1  },
'{ pfvf_port:1262  , pf:0 , vf:1262    , vf_active:1  },
'{ pfvf_port:1263  , pf:0 , vf:1263    , vf_active:1  },
'{ pfvf_port:1264  , pf:0 , vf:1264    , vf_active:1  },
'{ pfvf_port:1265  , pf:0 , vf:1265    , vf_active:1  },
'{ pfvf_port:1266  , pf:0 , vf:1266    , vf_active:1  },
'{ pfvf_port:1267  , pf:0 , vf:1267    , vf_active:1  },
'{ pfvf_port:1268  , pf:0 , vf:1268    , vf_active:1  },
'{ pfvf_port:1269  , pf:0 , vf:1269    , vf_active:1  },
'{ pfvf_port:1270  , pf:0 , vf:1270    , vf_active:1  },
'{ pfvf_port:1271  , pf:0 , vf:1271    , vf_active:1  },
'{ pfvf_port:1272  , pf:0 , vf:1272    , vf_active:1  },
'{ pfvf_port:1273  , pf:0 , vf:1273    , vf_active:1  },
'{ pfvf_port:1274  , pf:0 , vf:1274    , vf_active:1  },
'{ pfvf_port:1275  , pf:0 , vf:1275    , vf_active:1  },
'{ pfvf_port:1276  , pf:0 , vf:1276    , vf_active:1  },
'{ pfvf_port:1277  , pf:0 , vf:1277    , vf_active:1  },
'{ pfvf_port:1278  , pf:0 , vf:1278    , vf_active:1  },
'{ pfvf_port:1279  , pf:0 , vf:1279    , vf_active:1  },
'{ pfvf_port:1280  , pf:0 , vf:1280    , vf_active:1  },
'{ pfvf_port:1281  , pf:0 , vf:1281    , vf_active:1  },
'{ pfvf_port:1282  , pf:0 , vf:1282    , vf_active:1  },
'{ pfvf_port:1283  , pf:0 , vf:1283    , vf_active:1  },
'{ pfvf_port:1284  , pf:0 , vf:1284    , vf_active:1  },
'{ pfvf_port:1285  , pf:0 , vf:1285    , vf_active:1  },
'{ pfvf_port:1286  , pf:0 , vf:1286    , vf_active:1  },
'{ pfvf_port:1287  , pf:0 , vf:1287    , vf_active:1  },
'{ pfvf_port:1288  , pf:0 , vf:1288    , vf_active:1  },
'{ pfvf_port:1289  , pf:0 , vf:1289    , vf_active:1  },
'{ pfvf_port:1290  , pf:0 , vf:1290    , vf_active:1  },
'{ pfvf_port:1291  , pf:0 , vf:1291    , vf_active:1  },
'{ pfvf_port:1292  , pf:0 , vf:1292    , vf_active:1  },
'{ pfvf_port:1293  , pf:0 , vf:1293    , vf_active:1  },
'{ pfvf_port:1294  , pf:0 , vf:1294    , vf_active:1  },
'{ pfvf_port:1295  , pf:0 , vf:1295    , vf_active:1  },
'{ pfvf_port:1296  , pf:0 , vf:1296    , vf_active:1  },
'{ pfvf_port:1297  , pf:0 , vf:1297    , vf_active:1  },
'{ pfvf_port:1298  , pf:0 , vf:1298    , vf_active:1  },
'{ pfvf_port:1299  , pf:0 , vf:1299    , vf_active:1  },
'{ pfvf_port:1300  , pf:0 , vf:1300    , vf_active:1  },
'{ pfvf_port:1301  , pf:0 , vf:1301    , vf_active:1  },
'{ pfvf_port:1302  , pf:0 , vf:1302    , vf_active:1  },
'{ pfvf_port:1303  , pf:0 , vf:1303    , vf_active:1  },
'{ pfvf_port:1304  , pf:0 , vf:1304    , vf_active:1  },
'{ pfvf_port:1305  , pf:0 , vf:1305    , vf_active:1  },
'{ pfvf_port:1306  , pf:0 , vf:1306    , vf_active:1  },
'{ pfvf_port:1307  , pf:0 , vf:1307    , vf_active:1  },
'{ pfvf_port:1308  , pf:0 , vf:1308    , vf_active:1  },
'{ pfvf_port:1309  , pf:0 , vf:1309    , vf_active:1  },
'{ pfvf_port:1310  , pf:0 , vf:1310    , vf_active:1  },
'{ pfvf_port:1311  , pf:0 , vf:1311    , vf_active:1  },
'{ pfvf_port:1312  , pf:0 , vf:1312    , vf_active:1  },
'{ pfvf_port:1313  , pf:0 , vf:1313    , vf_active:1  },
'{ pfvf_port:1314  , pf:0 , vf:1314    , vf_active:1  },
'{ pfvf_port:1315  , pf:0 , vf:1315    , vf_active:1  },
'{ pfvf_port:1316  , pf:0 , vf:1316    , vf_active:1  },
'{ pfvf_port:1317  , pf:0 , vf:1317    , vf_active:1  },
'{ pfvf_port:1318  , pf:0 , vf:1318    , vf_active:1  },
'{ pfvf_port:1319  , pf:0 , vf:1319    , vf_active:1  },
'{ pfvf_port:1320  , pf:0 , vf:1320    , vf_active:1  },
'{ pfvf_port:1321  , pf:0 , vf:1321    , vf_active:1  },
'{ pfvf_port:1322  , pf:0 , vf:1322    , vf_active:1  },
'{ pfvf_port:1323  , pf:0 , vf:1323    , vf_active:1  },
'{ pfvf_port:1324  , pf:0 , vf:1324    , vf_active:1  },
'{ pfvf_port:1325  , pf:0 , vf:1325    , vf_active:1  },
'{ pfvf_port:1326  , pf:0 , vf:1326    , vf_active:1  },
'{ pfvf_port:1327  , pf:0 , vf:1327    , vf_active:1  },
'{ pfvf_port:1328  , pf:0 , vf:1328    , vf_active:1  },
'{ pfvf_port:1329  , pf:0 , vf:1329    , vf_active:1  },
'{ pfvf_port:1330  , pf:0 , vf:1330    , vf_active:1  },
'{ pfvf_port:1331  , pf:0 , vf:1331    , vf_active:1  },
'{ pfvf_port:1332  , pf:0 , vf:1332    , vf_active:1  },
'{ pfvf_port:1333  , pf:0 , vf:1333    , vf_active:1  },
'{ pfvf_port:1334  , pf:0 , vf:1334    , vf_active:1  },
'{ pfvf_port:1335  , pf:0 , vf:1335    , vf_active:1  },
'{ pfvf_port:1336  , pf:0 , vf:1336    , vf_active:1  },
'{ pfvf_port:1337  , pf:0 , vf:1337    , vf_active:1  },
'{ pfvf_port:1338  , pf:0 , vf:1338    , vf_active:1  },
'{ pfvf_port:1339  , pf:0 , vf:1339    , vf_active:1  },
'{ pfvf_port:1340  , pf:0 , vf:1340    , vf_active:1  },
'{ pfvf_port:1341  , pf:0 , vf:1341    , vf_active:1  },
'{ pfvf_port:1342  , pf:0 , vf:1342    , vf_active:1  },
'{ pfvf_port:1343  , pf:0 , vf:1343    , vf_active:1  },
'{ pfvf_port:1344  , pf:0 , vf:1344    , vf_active:1  },
'{ pfvf_port:1345  , pf:0 , vf:1345    , vf_active:1  },
'{ pfvf_port:1346  , pf:0 , vf:1346    , vf_active:1  },
'{ pfvf_port:1347  , pf:0 , vf:1347    , vf_active:1  },
'{ pfvf_port:1348  , pf:0 , vf:1348    , vf_active:1  },
'{ pfvf_port:1349  , pf:0 , vf:1349    , vf_active:1  },
'{ pfvf_port:1350  , pf:0 , vf:1350    , vf_active:1  },
'{ pfvf_port:1351  , pf:0 , vf:1351    , vf_active:1  },
'{ pfvf_port:1352  , pf:0 , vf:1352    , vf_active:1  },
'{ pfvf_port:1353  , pf:0 , vf:1353    , vf_active:1  },
'{ pfvf_port:1354  , pf:0 , vf:1354    , vf_active:1  },
'{ pfvf_port:1355  , pf:0 , vf:1355    , vf_active:1  },
'{ pfvf_port:1356  , pf:0 , vf:1356    , vf_active:1  },
'{ pfvf_port:1357  , pf:0 , vf:1357    , vf_active:1  },
'{ pfvf_port:1358  , pf:0 , vf:1358    , vf_active:1  },
'{ pfvf_port:1359  , pf:0 , vf:1359    , vf_active:1  },
'{ pfvf_port:1360  , pf:0 , vf:1360    , vf_active:1  },
'{ pfvf_port:1361  , pf:0 , vf:1361    , vf_active:1  },
'{ pfvf_port:1362  , pf:0 , vf:1362    , vf_active:1  },
'{ pfvf_port:1363  , pf:0 , vf:1363    , vf_active:1  },
'{ pfvf_port:1364  , pf:0 , vf:1364    , vf_active:1  },
'{ pfvf_port:1365  , pf:0 , vf:1365    , vf_active:1  },
'{ pfvf_port:1366  , pf:0 , vf:1366    , vf_active:1  },
'{ pfvf_port:1367  , pf:0 , vf:1367    , vf_active:1  },
'{ pfvf_port:1368  , pf:0 , vf:1368    , vf_active:1  },
'{ pfvf_port:1369  , pf:0 , vf:1369    , vf_active:1  },
'{ pfvf_port:1370  , pf:0 , vf:1370    , vf_active:1  },
'{ pfvf_port:1371  , pf:0 , vf:1371    , vf_active:1  },
'{ pfvf_port:1372  , pf:0 , vf:1372    , vf_active:1  },
'{ pfvf_port:1373  , pf:0 , vf:1373    , vf_active:1  },
'{ pfvf_port:1374  , pf:0 , vf:1374    , vf_active:1  },
'{ pfvf_port:1375  , pf:0 , vf:1375    , vf_active:1  },
'{ pfvf_port:1376  , pf:0 , vf:1376    , vf_active:1  },
'{ pfvf_port:1377  , pf:0 , vf:1377    , vf_active:1  },
'{ pfvf_port:1378  , pf:0 , vf:1378    , vf_active:1  },
'{ pfvf_port:1379  , pf:0 , vf:1379    , vf_active:1  },
'{ pfvf_port:1380  , pf:0 , vf:1380    , vf_active:1  },
'{ pfvf_port:1381  , pf:0 , vf:1381    , vf_active:1  },
'{ pfvf_port:1382  , pf:0 , vf:1382    , vf_active:1  },
'{ pfvf_port:1383  , pf:0 , vf:1383    , vf_active:1  },
'{ pfvf_port:1384  , pf:0 , vf:1384    , vf_active:1  },
'{ pfvf_port:1385  , pf:0 , vf:1385    , vf_active:1  },
'{ pfvf_port:1386  , pf:0 , vf:1386    , vf_active:1  },
'{ pfvf_port:1387  , pf:0 , vf:1387    , vf_active:1  },
'{ pfvf_port:1388  , pf:0 , vf:1388    , vf_active:1  },
'{ pfvf_port:1389  , pf:0 , vf:1389    , vf_active:1  },
'{ pfvf_port:1390  , pf:0 , vf:1390    , vf_active:1  },
'{ pfvf_port:1391  , pf:0 , vf:1391    , vf_active:1  },
'{ pfvf_port:1392  , pf:0 , vf:1392    , vf_active:1  },
'{ pfvf_port:1393  , pf:0 , vf:1393    , vf_active:1  },
'{ pfvf_port:1394  , pf:0 , vf:1394    , vf_active:1  },
'{ pfvf_port:1395  , pf:0 , vf:1395    , vf_active:1  },
'{ pfvf_port:1396  , pf:0 , vf:1396    , vf_active:1  },
'{ pfvf_port:1397  , pf:0 , vf:1397    , vf_active:1  },
'{ pfvf_port:1398  , pf:0 , vf:1398    , vf_active:1  },
'{ pfvf_port:1399  , pf:0 , vf:1399    , vf_active:1  },
'{ pfvf_port:1400  , pf:0 , vf:1400    , vf_active:1  },
'{ pfvf_port:1401  , pf:0 , vf:1401    , vf_active:1  },
'{ pfvf_port:1402  , pf:0 , vf:1402    , vf_active:1  },
'{ pfvf_port:1403  , pf:0 , vf:1403    , vf_active:1  },
'{ pfvf_port:1404  , pf:0 , vf:1404    , vf_active:1  },
'{ pfvf_port:1405  , pf:0 , vf:1405    , vf_active:1  },
'{ pfvf_port:1406  , pf:0 , vf:1406    , vf_active:1  },
'{ pfvf_port:1407  , pf:0 , vf:1407    , vf_active:1  },
'{ pfvf_port:1408  , pf:0 , vf:1408    , vf_active:1  },
'{ pfvf_port:1409  , pf:0 , vf:1409    , vf_active:1  },
'{ pfvf_port:1410  , pf:0 , vf:1410    , vf_active:1  },
'{ pfvf_port:1411  , pf:0 , vf:1411    , vf_active:1  },
'{ pfvf_port:1412  , pf:0 , vf:1412    , vf_active:1  },
'{ pfvf_port:1413  , pf:0 , vf:1413    , vf_active:1  },
'{ pfvf_port:1414  , pf:0 , vf:1414    , vf_active:1  },
'{ pfvf_port:1415  , pf:0 , vf:1415    , vf_active:1  },
'{ pfvf_port:1416  , pf:0 , vf:1416    , vf_active:1  },
'{ pfvf_port:1417  , pf:0 , vf:1417    , vf_active:1  },
'{ pfvf_port:1418  , pf:0 , vf:1418    , vf_active:1  },
'{ pfvf_port:1419  , pf:0 , vf:1419    , vf_active:1  },
'{ pfvf_port:1420  , pf:0 , vf:1420    , vf_active:1  },
'{ pfvf_port:1421  , pf:0 , vf:1421    , vf_active:1  },
'{ pfvf_port:1422  , pf:0 , vf:1422    , vf_active:1  },
'{ pfvf_port:1423  , pf:0 , vf:1423    , vf_active:1  },
'{ pfvf_port:1424  , pf:0 , vf:1424    , vf_active:1  },
'{ pfvf_port:1425  , pf:0 , vf:1425    , vf_active:1  },
'{ pfvf_port:1426  , pf:0 , vf:1426    , vf_active:1  },
'{ pfvf_port:1427  , pf:0 , vf:1427    , vf_active:1  },
'{ pfvf_port:1428  , pf:0 , vf:1428    , vf_active:1  },
'{ pfvf_port:1429  , pf:0 , vf:1429    , vf_active:1  },
'{ pfvf_port:1430  , pf:0 , vf:1430    , vf_active:1  },
'{ pfvf_port:1431  , pf:0 , vf:1431    , vf_active:1  },
'{ pfvf_port:1432  , pf:0 , vf:1432    , vf_active:1  },
'{ pfvf_port:1433  , pf:0 , vf:1433    , vf_active:1  },
'{ pfvf_port:1434  , pf:0 , vf:1434    , vf_active:1  },
'{ pfvf_port:1435  , pf:0 , vf:1435    , vf_active:1  },
'{ pfvf_port:1436  , pf:0 , vf:1436    , vf_active:1  },
'{ pfvf_port:1437  , pf:0 , vf:1437    , vf_active:1  },
'{ pfvf_port:1438  , pf:0 , vf:1438    , vf_active:1  },
'{ pfvf_port:1439  , pf:0 , vf:1439    , vf_active:1  },
'{ pfvf_port:1440  , pf:0 , vf:1440    , vf_active:1  },
'{ pfvf_port:1441  , pf:0 , vf:1441    , vf_active:1  },
'{ pfvf_port:1442  , pf:0 , vf:1442    , vf_active:1  },
'{ pfvf_port:1443  , pf:0 , vf:1443    , vf_active:1  },
'{ pfvf_port:1444  , pf:0 , vf:1444    , vf_active:1  },
'{ pfvf_port:1445  , pf:0 , vf:1445    , vf_active:1  },
'{ pfvf_port:1446  , pf:0 , vf:1446    , vf_active:1  },
'{ pfvf_port:1447  , pf:0 , vf:1447    , vf_active:1  },
'{ pfvf_port:1448  , pf:0 , vf:1448    , vf_active:1  },
'{ pfvf_port:1449  , pf:0 , vf:1449    , vf_active:1  },
'{ pfvf_port:1450  , pf:0 , vf:1450    , vf_active:1  },
'{ pfvf_port:1451  , pf:0 , vf:1451    , vf_active:1  },
'{ pfvf_port:1452  , pf:0 , vf:1452    , vf_active:1  },
'{ pfvf_port:1453  , pf:0 , vf:1453    , vf_active:1  },
'{ pfvf_port:1454  , pf:0 , vf:1454    , vf_active:1  },
'{ pfvf_port:1455  , pf:0 , vf:1455    , vf_active:1  },
'{ pfvf_port:1456  , pf:0 , vf:1456    , vf_active:1  },
'{ pfvf_port:1457  , pf:0 , vf:1457    , vf_active:1  },
'{ pfvf_port:1458  , pf:0 , vf:1458    , vf_active:1  },
'{ pfvf_port:1459  , pf:0 , vf:1459    , vf_active:1  },
'{ pfvf_port:1460  , pf:0 , vf:1460    , vf_active:1  },
'{ pfvf_port:1461  , pf:0 , vf:1461    , vf_active:1  },
'{ pfvf_port:1462  , pf:0 , vf:1462    , vf_active:1  },
'{ pfvf_port:1463  , pf:0 , vf:1463    , vf_active:1  },
'{ pfvf_port:1464  , pf:0 , vf:1464    , vf_active:1  },
'{ pfvf_port:1465  , pf:0 , vf:1465    , vf_active:1  },
'{ pfvf_port:1466  , pf:0 , vf:1466    , vf_active:1  },
'{ pfvf_port:1467  , pf:0 , vf:1467    , vf_active:1  },
'{ pfvf_port:1468  , pf:0 , vf:1468    , vf_active:1  },
'{ pfvf_port:1469  , pf:0 , vf:1469    , vf_active:1  },
'{ pfvf_port:1470  , pf:0 , vf:1470    , vf_active:1  },
'{ pfvf_port:1471  , pf:0 , vf:1471    , vf_active:1  },
'{ pfvf_port:1472  , pf:0 , vf:1472    , vf_active:1  },
'{ pfvf_port:1473  , pf:0 , vf:1473    , vf_active:1  },
'{ pfvf_port:1474  , pf:0 , vf:1474    , vf_active:1  },
'{ pfvf_port:1475  , pf:0 , vf:1475    , vf_active:1  },
'{ pfvf_port:1476  , pf:0 , vf:1476    , vf_active:1  },
'{ pfvf_port:1477  , pf:0 , vf:1477    , vf_active:1  },
'{ pfvf_port:1478  , pf:0 , vf:1478    , vf_active:1  },
'{ pfvf_port:1479  , pf:0 , vf:1479    , vf_active:1  },
'{ pfvf_port:1480  , pf:0 , vf:1480    , vf_active:1  },
'{ pfvf_port:1481  , pf:0 , vf:1481    , vf_active:1  },
'{ pfvf_port:1482  , pf:0 , vf:1482    , vf_active:1  },
'{ pfvf_port:1483  , pf:0 , vf:1483    , vf_active:1  },
'{ pfvf_port:1484  , pf:0 , vf:1484    , vf_active:1  },
'{ pfvf_port:1485  , pf:0 , vf:1485    , vf_active:1  },
'{ pfvf_port:1486  , pf:0 , vf:1486    , vf_active:1  },
'{ pfvf_port:1487  , pf:0 , vf:1487    , vf_active:1  },
'{ pfvf_port:1488  , pf:0 , vf:1488    , vf_active:1  },
'{ pfvf_port:1489  , pf:0 , vf:1489    , vf_active:1  },
'{ pfvf_port:1490  , pf:0 , vf:1490    , vf_active:1  },
'{ pfvf_port:1491  , pf:0 , vf:1491    , vf_active:1  },
'{ pfvf_port:1492  , pf:0 , vf:1492    , vf_active:1  },
'{ pfvf_port:1493  , pf:0 , vf:1493    , vf_active:1  },
'{ pfvf_port:1494  , pf:0 , vf:1494    , vf_active:1  },
'{ pfvf_port:1495  , pf:0 , vf:1495    , vf_active:1  },
'{ pfvf_port:1496  , pf:0 , vf:1496    , vf_active:1  },
'{ pfvf_port:1497  , pf:0 , vf:1497    , vf_active:1  },
'{ pfvf_port:1498  , pf:0 , vf:1498    , vf_active:1  },
'{ pfvf_port:1499  , pf:0 , vf:1499    , vf_active:1  },
'{ pfvf_port:1500  , pf:0 , vf:1500    , vf_active:1  },
'{ pfvf_port:1501  , pf:0 , vf:1501    , vf_active:1  },
'{ pfvf_port:1502  , pf:0 , vf:1502    , vf_active:1  },
'{ pfvf_port:1503  , pf:0 , vf:1503    , vf_active:1  },
'{ pfvf_port:1504  , pf:0 , vf:1504    , vf_active:1  },
'{ pfvf_port:1505  , pf:0 , vf:1505    , vf_active:1  },
'{ pfvf_port:1506  , pf:0 , vf:1506    , vf_active:1  },
'{ pfvf_port:1507  , pf:0 , vf:1507    , vf_active:1  },
'{ pfvf_port:1508  , pf:0 , vf:1508    , vf_active:1  },
'{ pfvf_port:1509  , pf:0 , vf:1509    , vf_active:1  },
'{ pfvf_port:1510  , pf:0 , vf:1510    , vf_active:1  },
'{ pfvf_port:1511  , pf:0 , vf:1511    , vf_active:1  },
'{ pfvf_port:1512  , pf:0 , vf:1512    , vf_active:1  },
'{ pfvf_port:1513  , pf:0 , vf:1513    , vf_active:1  },
'{ pfvf_port:1514  , pf:0 , vf:1514    , vf_active:1  },
'{ pfvf_port:1515  , pf:0 , vf:1515    , vf_active:1  },
'{ pfvf_port:1516  , pf:0 , vf:1516    , vf_active:1  },
'{ pfvf_port:1517  , pf:0 , vf:1517    , vf_active:1  },
'{ pfvf_port:1518  , pf:0 , vf:1518    , vf_active:1  },
'{ pfvf_port:1519  , pf:0 , vf:1519    , vf_active:1  },
'{ pfvf_port:1520  , pf:0 , vf:1520    , vf_active:1  },
'{ pfvf_port:1521  , pf:0 , vf:1521    , vf_active:1  },
'{ pfvf_port:1522  , pf:0 , vf:1522    , vf_active:1  },
'{ pfvf_port:1523  , pf:0 , vf:1523    , vf_active:1  },
'{ pfvf_port:1524  , pf:0 , vf:1524    , vf_active:1  },
'{ pfvf_port:1525  , pf:0 , vf:1525    , vf_active:1  },
'{ pfvf_port:1526  , pf:0 , vf:1526    , vf_active:1  },
'{ pfvf_port:1527  , pf:0 , vf:1527    , vf_active:1  },
'{ pfvf_port:1528  , pf:0 , vf:1528    , vf_active:1  },
'{ pfvf_port:1529  , pf:0 , vf:1529    , vf_active:1  },
'{ pfvf_port:1530  , pf:0 , vf:1530    , vf_active:1  },
'{ pfvf_port:1531  , pf:0 , vf:1531    , vf_active:1  },
'{ pfvf_port:1532  , pf:0 , vf:1532    , vf_active:1  },
'{ pfvf_port:1533  , pf:0 , vf:1533    , vf_active:1  },
'{ pfvf_port:1534  , pf:0 , vf:1534    , vf_active:1  },
'{ pfvf_port:1535  , pf:0 , vf:1535    , vf_active:1  },
'{ pfvf_port:1536  , pf:0 , vf:1536    , vf_active:1  },
'{ pfvf_port:1537  , pf:0 , vf:1537    , vf_active:1  },
'{ pfvf_port:1538  , pf:0 , vf:1538    , vf_active:1  },
'{ pfvf_port:1539  , pf:0 , vf:1539    , vf_active:1  },
'{ pfvf_port:1540  , pf:0 , vf:1540    , vf_active:1  },
'{ pfvf_port:1541  , pf:0 , vf:1541    , vf_active:1  },
'{ pfvf_port:1542  , pf:0 , vf:1542    , vf_active:1  },
'{ pfvf_port:1543  , pf:0 , vf:1543    , vf_active:1  },
'{ pfvf_port:1544  , pf:0 , vf:1544    , vf_active:1  },
'{ pfvf_port:1545  , pf:0 , vf:1545    , vf_active:1  },
'{ pfvf_port:1546  , pf:0 , vf:1546    , vf_active:1  },
'{ pfvf_port:1547  , pf:0 , vf:1547    , vf_active:1  },
'{ pfvf_port:1548  , pf:0 , vf:1548    , vf_active:1  },
'{ pfvf_port:1549  , pf:0 , vf:1549    , vf_active:1  },
'{ pfvf_port:1550  , pf:0 , vf:1550    , vf_active:1  },
'{ pfvf_port:1551  , pf:0 , vf:1551    , vf_active:1  },
'{ pfvf_port:1552  , pf:0 , vf:1552    , vf_active:1  },
'{ pfvf_port:1553  , pf:0 , vf:1553    , vf_active:1  },
'{ pfvf_port:1554  , pf:0 , vf:1554    , vf_active:1  },
'{ pfvf_port:1555  , pf:0 , vf:1555    , vf_active:1  },
'{ pfvf_port:1556  , pf:0 , vf:1556    , vf_active:1  },
'{ pfvf_port:1557  , pf:0 , vf:1557    , vf_active:1  },
'{ pfvf_port:1558  , pf:0 , vf:1558    , vf_active:1  },
'{ pfvf_port:1559  , pf:0 , vf:1559    , vf_active:1  },
'{ pfvf_port:1560  , pf:0 , vf:1560    , vf_active:1  },
'{ pfvf_port:1561  , pf:0 , vf:1561    , vf_active:1  },
'{ pfvf_port:1562  , pf:0 , vf:1562    , vf_active:1  },
'{ pfvf_port:1563  , pf:0 , vf:1563    , vf_active:1  },
'{ pfvf_port:1564  , pf:0 , vf:1564    , vf_active:1  },
'{ pfvf_port:1565  , pf:0 , vf:1565    , vf_active:1  },
'{ pfvf_port:1566  , pf:0 , vf:1566    , vf_active:1  },
'{ pfvf_port:1567  , pf:0 , vf:1567    , vf_active:1  },
'{ pfvf_port:1568  , pf:0 , vf:1568    , vf_active:1  },
'{ pfvf_port:1569  , pf:0 , vf:1569    , vf_active:1  },
'{ pfvf_port:1570  , pf:0 , vf:1570    , vf_active:1  },
'{ pfvf_port:1571  , pf:0 , vf:1571    , vf_active:1  },
'{ pfvf_port:1572  , pf:0 , vf:1572    , vf_active:1  },
'{ pfvf_port:1573  , pf:0 , vf:1573    , vf_active:1  },
'{ pfvf_port:1574  , pf:0 , vf:1574    , vf_active:1  },
'{ pfvf_port:1575  , pf:0 , vf:1575    , vf_active:1  },
'{ pfvf_port:1576  , pf:0 , vf:1576    , vf_active:1  },
'{ pfvf_port:1577  , pf:0 , vf:1577    , vf_active:1  },
'{ pfvf_port:1578  , pf:0 , vf:1578    , vf_active:1  },
'{ pfvf_port:1579  , pf:0 , vf:1579    , vf_active:1  },
'{ pfvf_port:1580  , pf:0 , vf:1580    , vf_active:1  },
'{ pfvf_port:1581  , pf:0 , vf:1581    , vf_active:1  },
'{ pfvf_port:1582  , pf:0 , vf:1582    , vf_active:1  },
'{ pfvf_port:1583  , pf:0 , vf:1583    , vf_active:1  },
'{ pfvf_port:1584  , pf:0 , vf:1584    , vf_active:1  },
'{ pfvf_port:1585  , pf:0 , vf:1585    , vf_active:1  },
'{ pfvf_port:1586  , pf:0 , vf:1586    , vf_active:1  },
'{ pfvf_port:1587  , pf:0 , vf:1587    , vf_active:1  },
'{ pfvf_port:1588  , pf:0 , vf:1588    , vf_active:1  },
'{ pfvf_port:1589  , pf:0 , vf:1589    , vf_active:1  },
'{ pfvf_port:1590  , pf:0 , vf:1590    , vf_active:1  },
'{ pfvf_port:1591  , pf:0 , vf:1591    , vf_active:1  },
'{ pfvf_port:1592  , pf:0 , vf:1592    , vf_active:1  },
'{ pfvf_port:1593  , pf:0 , vf:1593    , vf_active:1  },
'{ pfvf_port:1594  , pf:0 , vf:1594    , vf_active:1  },
'{ pfvf_port:1595  , pf:0 , vf:1595    , vf_active:1  },
'{ pfvf_port:1596  , pf:0 , vf:1596    , vf_active:1  },
'{ pfvf_port:1597  , pf:0 , vf:1597    , vf_active:1  },
'{ pfvf_port:1598  , pf:0 , vf:1598    , vf_active:1  },
'{ pfvf_port:1599  , pf:0 , vf:1599    , vf_active:1  },
'{ pfvf_port:1600  , pf:0 , vf:1600    , vf_active:1  },
'{ pfvf_port:1601  , pf:0 , vf:1601    , vf_active:1  },
'{ pfvf_port:1602  , pf:0 , vf:1602    , vf_active:1  },
'{ pfvf_port:1603  , pf:0 , vf:1603    , vf_active:1  },
'{ pfvf_port:1604  , pf:0 , vf:1604    , vf_active:1  },
'{ pfvf_port:1605  , pf:0 , vf:1605    , vf_active:1  },
'{ pfvf_port:1606  , pf:0 , vf:1606    , vf_active:1  },
'{ pfvf_port:1607  , pf:0 , vf:1607    , vf_active:1  },
'{ pfvf_port:1608  , pf:0 , vf:1608    , vf_active:1  },
'{ pfvf_port:1609  , pf:0 , vf:1609    , vf_active:1  },
'{ pfvf_port:1610  , pf:0 , vf:1610    , vf_active:1  },
'{ pfvf_port:1611  , pf:0 , vf:1611    , vf_active:1  },
'{ pfvf_port:1612  , pf:0 , vf:1612    , vf_active:1  },
'{ pfvf_port:1613  , pf:0 , vf:1613    , vf_active:1  },
'{ pfvf_port:1614  , pf:0 , vf:1614    , vf_active:1  },
'{ pfvf_port:1615  , pf:0 , vf:1615    , vf_active:1  },
'{ pfvf_port:1616  , pf:0 , vf:1616    , vf_active:1  },
'{ pfvf_port:1617  , pf:0 , vf:1617    , vf_active:1  },
'{ pfvf_port:1618  , pf:0 , vf:1618    , vf_active:1  },
'{ pfvf_port:1619  , pf:0 , vf:1619    , vf_active:1  },
'{ pfvf_port:1620  , pf:0 , vf:1620    , vf_active:1  },
'{ pfvf_port:1621  , pf:0 , vf:1621    , vf_active:1  },
'{ pfvf_port:1622  , pf:0 , vf:1622    , vf_active:1  },
'{ pfvf_port:1623  , pf:0 , vf:1623    , vf_active:1  },
'{ pfvf_port:1624  , pf:0 , vf:1624    , vf_active:1  },
'{ pfvf_port:1625  , pf:0 , vf:1625    , vf_active:1  },
'{ pfvf_port:1626  , pf:0 , vf:1626    , vf_active:1  },
'{ pfvf_port:1627  , pf:0 , vf:1627    , vf_active:1  },
'{ pfvf_port:1628  , pf:0 , vf:1628    , vf_active:1  },
'{ pfvf_port:1629  , pf:0 , vf:1629    , vf_active:1  },
'{ pfvf_port:1630  , pf:0 , vf:1630    , vf_active:1  },
'{ pfvf_port:1631  , pf:0 , vf:1631    , vf_active:1  },
'{ pfvf_port:1632  , pf:0 , vf:1632    , vf_active:1  },
'{ pfvf_port:1633  , pf:0 , vf:1633    , vf_active:1  },
'{ pfvf_port:1634  , pf:0 , vf:1634    , vf_active:1  },
'{ pfvf_port:1635  , pf:0 , vf:1635    , vf_active:1  },
'{ pfvf_port:1636  , pf:0 , vf:1636    , vf_active:1  },
'{ pfvf_port:1637  , pf:0 , vf:1637    , vf_active:1  },
'{ pfvf_port:1638  , pf:0 , vf:1638    , vf_active:1  },
'{ pfvf_port:1639  , pf:0 , vf:1639    , vf_active:1  },
'{ pfvf_port:1640  , pf:0 , vf:1640    , vf_active:1  },
'{ pfvf_port:1641  , pf:0 , vf:1641    , vf_active:1  },
'{ pfvf_port:1642  , pf:0 , vf:1642    , vf_active:1  },
'{ pfvf_port:1643  , pf:0 , vf:1643    , vf_active:1  },
'{ pfvf_port:1644  , pf:0 , vf:1644    , vf_active:1  },
'{ pfvf_port:1645  , pf:0 , vf:1645    , vf_active:1  },
'{ pfvf_port:1646  , pf:0 , vf:1646    , vf_active:1  },
'{ pfvf_port:1647  , pf:0 , vf:1647    , vf_active:1  },
'{ pfvf_port:1648  , pf:0 , vf:1648    , vf_active:1  },
'{ pfvf_port:1649  , pf:0 , vf:1649    , vf_active:1  },
'{ pfvf_port:1650  , pf:0 , vf:1650    , vf_active:1  },
'{ pfvf_port:1651  , pf:0 , vf:1651    , vf_active:1  },
'{ pfvf_port:1652  , pf:0 , vf:1652    , vf_active:1  },
'{ pfvf_port:1653  , pf:0 , vf:1653    , vf_active:1  },
'{ pfvf_port:1654  , pf:0 , vf:1654    , vf_active:1  },
'{ pfvf_port:1655  , pf:0 , vf:1655    , vf_active:1  },
'{ pfvf_port:1656  , pf:0 , vf:1656    , vf_active:1  },
'{ pfvf_port:1657  , pf:0 , vf:1657    , vf_active:1  },
'{ pfvf_port:1658  , pf:0 , vf:1658    , vf_active:1  },
'{ pfvf_port:1659  , pf:0 , vf:1659    , vf_active:1  },
'{ pfvf_port:1660  , pf:0 , vf:1660    , vf_active:1  },
'{ pfvf_port:1661  , pf:0 , vf:1661    , vf_active:1  },
'{ pfvf_port:1662  , pf:0 , vf:1662    , vf_active:1  },
'{ pfvf_port:1663  , pf:0 , vf:1663    , vf_active:1  },
'{ pfvf_port:1664  , pf:0 , vf:1664    , vf_active:1  },
'{ pfvf_port:1665  , pf:0 , vf:1665    , vf_active:1  },
'{ pfvf_port:1666  , pf:0 , vf:1666    , vf_active:1  },
'{ pfvf_port:1667  , pf:0 , vf:1667    , vf_active:1  },
'{ pfvf_port:1668  , pf:0 , vf:1668    , vf_active:1  },
'{ pfvf_port:1669  , pf:0 , vf:1669    , vf_active:1  },
'{ pfvf_port:1670  , pf:0 , vf:1670    , vf_active:1  },
'{ pfvf_port:1671  , pf:0 , vf:1671    , vf_active:1  },
'{ pfvf_port:1672  , pf:0 , vf:1672    , vf_active:1  },
'{ pfvf_port:1673  , pf:0 , vf:1673    , vf_active:1  },
'{ pfvf_port:1674  , pf:0 , vf:1674    , vf_active:1  },
'{ pfvf_port:1675  , pf:0 , vf:1675    , vf_active:1  },
'{ pfvf_port:1676  , pf:0 , vf:1676    , vf_active:1  },
'{ pfvf_port:1677  , pf:0 , vf:1677    , vf_active:1  },
'{ pfvf_port:1678  , pf:0 , vf:1678    , vf_active:1  },
'{ pfvf_port:1679  , pf:0 , vf:1679    , vf_active:1  },
'{ pfvf_port:1680  , pf:0 , vf:1680    , vf_active:1  },
'{ pfvf_port:1681  , pf:0 , vf:1681    , vf_active:1  },
'{ pfvf_port:1682  , pf:0 , vf:1682    , vf_active:1  },
'{ pfvf_port:1683  , pf:0 , vf:1683    , vf_active:1  },
'{ pfvf_port:1684  , pf:0 , vf:1684    , vf_active:1  },
'{ pfvf_port:1685  , pf:0 , vf:1685    , vf_active:1  },
'{ pfvf_port:1686  , pf:0 , vf:1686    , vf_active:1  },
'{ pfvf_port:1687  , pf:0 , vf:1687    , vf_active:1  },
'{ pfvf_port:1688  , pf:0 , vf:1688    , vf_active:1  },
'{ pfvf_port:1689  , pf:0 , vf:1689    , vf_active:1  },
'{ pfvf_port:1690  , pf:0 , vf:1690    , vf_active:1  },
'{ pfvf_port:1691  , pf:0 , vf:1691    , vf_active:1  },
'{ pfvf_port:1692  , pf:0 , vf:1692    , vf_active:1  },
'{ pfvf_port:1693  , pf:0 , vf:1693    , vf_active:1  },
'{ pfvf_port:1694  , pf:0 , vf:1694    , vf_active:1  },
'{ pfvf_port:1695  , pf:0 , vf:1695    , vf_active:1  },
'{ pfvf_port:1696  , pf:0 , vf:1696    , vf_active:1  },
'{ pfvf_port:1697  , pf:0 , vf:1697    , vf_active:1  },
'{ pfvf_port:1698  , pf:0 , vf:1698    , vf_active:1  },
'{ pfvf_port:1699  , pf:0 , vf:1699    , vf_active:1  },
'{ pfvf_port:1700  , pf:0 , vf:1700    , vf_active:1  },
'{ pfvf_port:1701  , pf:0 , vf:1701    , vf_active:1  },
'{ pfvf_port:1702  , pf:0 , vf:1702    , vf_active:1  },
'{ pfvf_port:1703  , pf:0 , vf:1703    , vf_active:1  },
'{ pfvf_port:1704  , pf:0 , vf:1704    , vf_active:1  },
'{ pfvf_port:1705  , pf:0 , vf:1705    , vf_active:1  },
'{ pfvf_port:1706  , pf:0 , vf:1706    , vf_active:1  },
'{ pfvf_port:1707  , pf:0 , vf:1707    , vf_active:1  },
'{ pfvf_port:1708  , pf:0 , vf:1708    , vf_active:1  },
'{ pfvf_port:1709  , pf:0 , vf:1709    , vf_active:1  },
'{ pfvf_port:1710  , pf:0 , vf:1710    , vf_active:1  },
'{ pfvf_port:1711  , pf:0 , vf:1711    , vf_active:1  },
'{ pfvf_port:1712  , pf:0 , vf:1712    , vf_active:1  },
'{ pfvf_port:1713  , pf:0 , vf:1713    , vf_active:1  },
'{ pfvf_port:1714  , pf:0 , vf:1714    , vf_active:1  },
'{ pfvf_port:1715  , pf:0 , vf:1715    , vf_active:1  },
'{ pfvf_port:1716  , pf:0 , vf:1716    , vf_active:1  },
'{ pfvf_port:1717  , pf:0 , vf:1717    , vf_active:1  },
'{ pfvf_port:1718  , pf:0 , vf:1718    , vf_active:1  },
'{ pfvf_port:1719  , pf:0 , vf:1719    , vf_active:1  },
'{ pfvf_port:1720  , pf:0 , vf:1720    , vf_active:1  },
'{ pfvf_port:1721  , pf:0 , vf:1721    , vf_active:1  },
'{ pfvf_port:1722  , pf:0 , vf:1722    , vf_active:1  },
'{ pfvf_port:1723  , pf:0 , vf:1723    , vf_active:1  },
'{ pfvf_port:1724  , pf:0 , vf:1724    , vf_active:1  },
'{ pfvf_port:1725  , pf:0 , vf:1725    , vf_active:1  },
'{ pfvf_port:1726  , pf:0 , vf:1726    , vf_active:1  },
'{ pfvf_port:1727  , pf:0 , vf:1727    , vf_active:1  },
'{ pfvf_port:1728  , pf:0 , vf:1728    , vf_active:1  },
'{ pfvf_port:1729  , pf:0 , vf:1729    , vf_active:1  },
'{ pfvf_port:1730  , pf:0 , vf:1730    , vf_active:1  },
'{ pfvf_port:1731  , pf:0 , vf:1731    , vf_active:1  },
'{ pfvf_port:1732  , pf:0 , vf:1732    , vf_active:1  },
'{ pfvf_port:1733  , pf:0 , vf:1733    , vf_active:1  },
'{ pfvf_port:1734  , pf:0 , vf:1734    , vf_active:1  },
'{ pfvf_port:1735  , pf:0 , vf:1735    , vf_active:1  },
'{ pfvf_port:1736  , pf:0 , vf:1736    , vf_active:1  },
'{ pfvf_port:1737  , pf:0 , vf:1737    , vf_active:1  },
'{ pfvf_port:1738  , pf:0 , vf:1738    , vf_active:1  },
'{ pfvf_port:1739  , pf:0 , vf:1739    , vf_active:1  },
'{ pfvf_port:1740  , pf:0 , vf:1740    , vf_active:1  },
'{ pfvf_port:1741  , pf:0 , vf:1741    , vf_active:1  },
'{ pfvf_port:1742  , pf:0 , vf:1742    , vf_active:1  },
'{ pfvf_port:1743  , pf:0 , vf:1743    , vf_active:1  },
'{ pfvf_port:1744  , pf:0 , vf:1744    , vf_active:1  },
'{ pfvf_port:1745  , pf:0 , vf:1745    , vf_active:1  },
'{ pfvf_port:1746  , pf:0 , vf:1746    , vf_active:1  },
'{ pfvf_port:1747  , pf:0 , vf:1747    , vf_active:1  },
'{ pfvf_port:1748  , pf:0 , vf:1748    , vf_active:1  },
'{ pfvf_port:1749  , pf:0 , vf:1749    , vf_active:1  },
'{ pfvf_port:1750  , pf:0 , vf:1750    , vf_active:1  },
'{ pfvf_port:1751  , pf:0 , vf:1751    , vf_active:1  },
'{ pfvf_port:1752  , pf:0 , vf:1752    , vf_active:1  },
'{ pfvf_port:1753  , pf:0 , vf:1753    , vf_active:1  },
'{ pfvf_port:1754  , pf:0 , vf:1754    , vf_active:1  },
'{ pfvf_port:1755  , pf:0 , vf:1755    , vf_active:1  },
'{ pfvf_port:1756  , pf:0 , vf:1756    , vf_active:1  },
'{ pfvf_port:1757  , pf:0 , vf:1757    , vf_active:1  },
'{ pfvf_port:1758  , pf:0 , vf:1758    , vf_active:1  },
'{ pfvf_port:1759  , pf:0 , vf:1759    , vf_active:1  },
'{ pfvf_port:1760  , pf:0 , vf:1760    , vf_active:1  },
'{ pfvf_port:1761  , pf:0 , vf:1761    , vf_active:1  },
'{ pfvf_port:1762  , pf:0 , vf:1762    , vf_active:1  },
'{ pfvf_port:1763  , pf:0 , vf:1763    , vf_active:1  },
'{ pfvf_port:1764  , pf:0 , vf:1764    , vf_active:1  },
'{ pfvf_port:1765  , pf:0 , vf:1765    , vf_active:1  },
'{ pfvf_port:1766  , pf:0 , vf:1766    , vf_active:1  },
'{ pfvf_port:1767  , pf:0 , vf:1767    , vf_active:1  },
'{ pfvf_port:1768  , pf:0 , vf:1768    , vf_active:1  },
'{ pfvf_port:1769  , pf:0 , vf:1769    , vf_active:1  },
'{ pfvf_port:1770  , pf:0 , vf:1770    , vf_active:1  },
'{ pfvf_port:1771  , pf:0 , vf:1771    , vf_active:1  },
'{ pfvf_port:1772  , pf:0 , vf:1772    , vf_active:1  },
'{ pfvf_port:1773  , pf:0 , vf:1773    , vf_active:1  },
'{ pfvf_port:1774  , pf:0 , vf:1774    , vf_active:1  },
'{ pfvf_port:1775  , pf:0 , vf:1775    , vf_active:1  },
'{ pfvf_port:1776  , pf:0 , vf:1776    , vf_active:1  },
'{ pfvf_port:1777  , pf:0 , vf:1777    , vf_active:1  },
'{ pfvf_port:1778  , pf:0 , vf:1778    , vf_active:1  },
'{ pfvf_port:1779  , pf:0 , vf:1779    , vf_active:1  },
'{ pfvf_port:1780  , pf:0 , vf:1780    , vf_active:1  },
'{ pfvf_port:1781  , pf:0 , vf:1781    , vf_active:1  },
'{ pfvf_port:1782  , pf:0 , vf:1782    , vf_active:1  },
'{ pfvf_port:1783  , pf:0 , vf:1783    , vf_active:1  },
'{ pfvf_port:1784  , pf:0 , vf:1784    , vf_active:1  },
'{ pfvf_port:1785  , pf:0 , vf:1785    , vf_active:1  },
'{ pfvf_port:1786  , pf:0 , vf:1786    , vf_active:1  },
'{ pfvf_port:1787  , pf:0 , vf:1787    , vf_active:1  },
'{ pfvf_port:1788  , pf:0 , vf:1788    , vf_active:1  },
'{ pfvf_port:1789  , pf:0 , vf:1789    , vf_active:1  },
'{ pfvf_port:1790  , pf:0 , vf:1790    , vf_active:1  },
'{ pfvf_port:1791  , pf:0 , vf:1791    , vf_active:1  },
'{ pfvf_port:1792  , pf:0 , vf:1792    , vf_active:1  },
'{ pfvf_port:1793  , pf:0 , vf:1793    , vf_active:1  },
'{ pfvf_port:1794  , pf:0 , vf:1794    , vf_active:1  },
'{ pfvf_port:1795  , pf:0 , vf:1795    , vf_active:1  },
'{ pfvf_port:1796  , pf:0 , vf:1796    , vf_active:1  },
'{ pfvf_port:1797  , pf:0 , vf:1797    , vf_active:1  },
'{ pfvf_port:1798  , pf:0 , vf:1798    , vf_active:1  },
'{ pfvf_port:1799  , pf:0 , vf:1799    , vf_active:1  },
'{ pfvf_port:1800  , pf:0 , vf:1800    , vf_active:1  },
'{ pfvf_port:1801  , pf:0 , vf:1801    , vf_active:1  },
'{ pfvf_port:1802  , pf:0 , vf:1802    , vf_active:1  },
'{ pfvf_port:1803  , pf:0 , vf:1803    , vf_active:1  },
'{ pfvf_port:1804  , pf:0 , vf:1804    , vf_active:1  },
'{ pfvf_port:1805  , pf:0 , vf:1805    , vf_active:1  },
'{ pfvf_port:1806  , pf:0 , vf:1806    , vf_active:1  },
'{ pfvf_port:1807  , pf:0 , vf:1807    , vf_active:1  },
'{ pfvf_port:1808  , pf:0 , vf:1808    , vf_active:1  },
'{ pfvf_port:1809  , pf:0 , vf:1809    , vf_active:1  },
'{ pfvf_port:1810  , pf:0 , vf:1810    , vf_active:1  },
'{ pfvf_port:1811  , pf:0 , vf:1811    , vf_active:1  },
'{ pfvf_port:1812  , pf:0 , vf:1812    , vf_active:1  },
'{ pfvf_port:1813  , pf:0 , vf:1813    , vf_active:1  },
'{ pfvf_port:1814  , pf:0 , vf:1814    , vf_active:1  },
'{ pfvf_port:1815  , pf:0 , vf:1815    , vf_active:1  },
'{ pfvf_port:1816  , pf:0 , vf:1816    , vf_active:1  },
'{ pfvf_port:1817  , pf:0 , vf:1817    , vf_active:1  },
'{ pfvf_port:1818  , pf:0 , vf:1818    , vf_active:1  },
'{ pfvf_port:1819  , pf:0 , vf:1819    , vf_active:1  },
'{ pfvf_port:1820  , pf:0 , vf:1820    , vf_active:1  },
'{ pfvf_port:1821  , pf:0 , vf:1821    , vf_active:1  },
'{ pfvf_port:1822  , pf:0 , vf:1822    , vf_active:1  },
'{ pfvf_port:1823  , pf:0 , vf:1823    , vf_active:1  },
'{ pfvf_port:1824  , pf:0 , vf:1824    , vf_active:1  },
'{ pfvf_port:1825  , pf:0 , vf:1825    , vf_active:1  },
'{ pfvf_port:1826  , pf:0 , vf:1826    , vf_active:1  },
'{ pfvf_port:1827  , pf:0 , vf:1827    , vf_active:1  },
'{ pfvf_port:1828  , pf:0 , vf:1828    , vf_active:1  },
'{ pfvf_port:1829  , pf:0 , vf:1829    , vf_active:1  },
'{ pfvf_port:1830  , pf:0 , vf:1830    , vf_active:1  },
'{ pfvf_port:1831  , pf:0 , vf:1831    , vf_active:1  },
'{ pfvf_port:1832  , pf:0 , vf:1832    , vf_active:1  },
'{ pfvf_port:1833  , pf:0 , vf:1833    , vf_active:1  },
'{ pfvf_port:1834  , pf:0 , vf:1834    , vf_active:1  },
'{ pfvf_port:1835  , pf:0 , vf:1835    , vf_active:1  },
'{ pfvf_port:1836  , pf:0 , vf:1836    , vf_active:1  },
'{ pfvf_port:1837  , pf:0 , vf:1837    , vf_active:1  },
'{ pfvf_port:1838  , pf:0 , vf:1838    , vf_active:1  },
'{ pfvf_port:1839  , pf:0 , vf:1839    , vf_active:1  },
'{ pfvf_port:1840  , pf:0 , vf:1840    , vf_active:1  },
'{ pfvf_port:1841  , pf:0 , vf:1841    , vf_active:1  },
'{ pfvf_port:1842  , pf:0 , vf:1842    , vf_active:1  },
'{ pfvf_port:1843  , pf:0 , vf:1843    , vf_active:1  },
'{ pfvf_port:1844  , pf:0 , vf:1844    , vf_active:1  },
'{ pfvf_port:1845  , pf:0 , vf:1845    , vf_active:1  },
'{ pfvf_port:1846  , pf:0 , vf:1846    , vf_active:1  },
'{ pfvf_port:1847  , pf:0 , vf:1847    , vf_active:1  },
'{ pfvf_port:1848  , pf:0 , vf:1848    , vf_active:1  },
'{ pfvf_port:1849  , pf:0 , vf:1849    , vf_active:1  },
'{ pfvf_port:1850  , pf:0 , vf:1850    , vf_active:1  },
'{ pfvf_port:1851  , pf:0 , vf:1851    , vf_active:1  },
'{ pfvf_port:1852  , pf:0 , vf:1852    , vf_active:1  },
'{ pfvf_port:1853  , pf:0 , vf:1853    , vf_active:1  },
'{ pfvf_port:1854  , pf:0 , vf:1854    , vf_active:1  },
'{ pfvf_port:1855  , pf:0 , vf:1855    , vf_active:1  },
'{ pfvf_port:1856  , pf:0 , vf:1856    , vf_active:1  },
'{ pfvf_port:1857  , pf:0 , vf:1857    , vf_active:1  },
'{ pfvf_port:1858  , pf:0 , vf:1858    , vf_active:1  },
'{ pfvf_port:1859  , pf:0 , vf:1859    , vf_active:1  },
'{ pfvf_port:1860  , pf:0 , vf:1860    , vf_active:1  },
'{ pfvf_port:1861  , pf:0 , vf:1861    , vf_active:1  },
'{ pfvf_port:1862  , pf:0 , vf:1862    , vf_active:1  },
'{ pfvf_port:1863  , pf:0 , vf:1863    , vf_active:1  },
'{ pfvf_port:1864  , pf:0 , vf:1864    , vf_active:1  },
'{ pfvf_port:1865  , pf:0 , vf:1865    , vf_active:1  },
'{ pfvf_port:1866  , pf:0 , vf:1866    , vf_active:1  },
'{ pfvf_port:1867  , pf:0 , vf:1867    , vf_active:1  },
'{ pfvf_port:1868  , pf:0 , vf:1868    , vf_active:1  },
'{ pfvf_port:1869  , pf:0 , vf:1869    , vf_active:1  },
'{ pfvf_port:1870  , pf:0 , vf:1870    , vf_active:1  },
'{ pfvf_port:1871  , pf:0 , vf:1871    , vf_active:1  },
'{ pfvf_port:1872  , pf:0 , vf:1872    , vf_active:1  },
'{ pfvf_port:1873  , pf:0 , vf:1873    , vf_active:1  },
'{ pfvf_port:1874  , pf:0 , vf:1874    , vf_active:1  },
'{ pfvf_port:1875  , pf:0 , vf:1875    , vf_active:1  },
'{ pfvf_port:1876  , pf:0 , vf:1876    , vf_active:1  },
'{ pfvf_port:1877  , pf:0 , vf:1877    , vf_active:1  },
'{ pfvf_port:1878  , pf:0 , vf:1878    , vf_active:1  },
'{ pfvf_port:1879  , pf:0 , vf:1879    , vf_active:1  },
'{ pfvf_port:1880  , pf:0 , vf:1880    , vf_active:1  },
'{ pfvf_port:1881  , pf:0 , vf:1881    , vf_active:1  },
'{ pfvf_port:1882  , pf:0 , vf:1882    , vf_active:1  },
'{ pfvf_port:1883  , pf:0 , vf:1883    , vf_active:1  },
'{ pfvf_port:1884  , pf:0 , vf:1884    , vf_active:1  },
'{ pfvf_port:1885  , pf:0 , vf:1885    , vf_active:1  },
'{ pfvf_port:1886  , pf:0 , vf:1886    , vf_active:1  },
'{ pfvf_port:1887  , pf:0 , vf:1887    , vf_active:1  },
'{ pfvf_port:1888  , pf:0 , vf:1888    , vf_active:1  },
'{ pfvf_port:1889  , pf:0 , vf:1889    , vf_active:1  },
'{ pfvf_port:1890  , pf:0 , vf:1890    , vf_active:1  },
'{ pfvf_port:1891  , pf:0 , vf:1891    , vf_active:1  },
'{ pfvf_port:1892  , pf:0 , vf:1892    , vf_active:1  },
'{ pfvf_port:1893  , pf:0 , vf:1893    , vf_active:1  },
'{ pfvf_port:1894  , pf:0 , vf:1894    , vf_active:1  },
'{ pfvf_port:1895  , pf:0 , vf:1895    , vf_active:1  },
'{ pfvf_port:1896  , pf:0 , vf:1896    , vf_active:1  },
'{ pfvf_port:1897  , pf:0 , vf:1897    , vf_active:1  },
'{ pfvf_port:1898  , pf:0 , vf:1898    , vf_active:1  },
'{ pfvf_port:1899  , pf:0 , vf:1899    , vf_active:1  },
'{ pfvf_port:1900  , pf:0 , vf:1900    , vf_active:1  },
'{ pfvf_port:1901  , pf:0 , vf:1901    , vf_active:1  },
'{ pfvf_port:1902  , pf:0 , vf:1902    , vf_active:1  },
'{ pfvf_port:1903  , pf:0 , vf:1903    , vf_active:1  },
'{ pfvf_port:1904  , pf:0 , vf:1904    , vf_active:1  },
'{ pfvf_port:1905  , pf:0 , vf:1905    , vf_active:1  },
'{ pfvf_port:1906  , pf:0 , vf:1906    , vf_active:1  },
'{ pfvf_port:1907  , pf:0 , vf:1907    , vf_active:1  },
'{ pfvf_port:1908  , pf:0 , vf:1908    , vf_active:1  },
'{ pfvf_port:1909  , pf:0 , vf:1909    , vf_active:1  },
'{ pfvf_port:1910  , pf:0 , vf:1910    , vf_active:1  },
'{ pfvf_port:1911  , pf:0 , vf:1911    , vf_active:1  },
'{ pfvf_port:1912  , pf:0 , vf:1912    , vf_active:1  },
'{ pfvf_port:1913  , pf:0 , vf:1913    , vf_active:1  },
'{ pfvf_port:1914  , pf:0 , vf:1914    , vf_active:1  },
'{ pfvf_port:1915  , pf:0 , vf:1915    , vf_active:1  },
'{ pfvf_port:1916  , pf:0 , vf:1916    , vf_active:1  },
'{ pfvf_port:1917  , pf:0 , vf:1917    , vf_active:1  },
'{ pfvf_port:1918  , pf:0 , vf:1918    , vf_active:1  },
'{ pfvf_port:1919  , pf:0 , vf:1919    , vf_active:1  },
'{ pfvf_port:1920  , pf:0 , vf:1920    , vf_active:1  },
'{ pfvf_port:1921  , pf:0 , vf:1921    , vf_active:1  },
'{ pfvf_port:1922  , pf:0 , vf:1922    , vf_active:1  },
'{ pfvf_port:1923  , pf:0 , vf:1923    , vf_active:1  },
'{ pfvf_port:1924  , pf:0 , vf:1924    , vf_active:1  },
'{ pfvf_port:1925  , pf:0 , vf:1925    , vf_active:1  },
'{ pfvf_port:1926  , pf:0 , vf:1926    , vf_active:1  },
'{ pfvf_port:1927  , pf:0 , vf:1927    , vf_active:1  },
'{ pfvf_port:1928  , pf:0 , vf:1928    , vf_active:1  },
'{ pfvf_port:1929  , pf:0 , vf:1929    , vf_active:1  },
'{ pfvf_port:1930  , pf:0 , vf:1930    , vf_active:1  },
'{ pfvf_port:1931  , pf:0 , vf:1931    , vf_active:1  },
'{ pfvf_port:1932  , pf:0 , vf:1932    , vf_active:1  },
'{ pfvf_port:1933  , pf:0 , vf:1933    , vf_active:1  },
'{ pfvf_port:1934  , pf:0 , vf:1934    , vf_active:1  },
'{ pfvf_port:1935  , pf:0 , vf:1935    , vf_active:1  },
'{ pfvf_port:1936  , pf:0 , vf:1936    , vf_active:1  },
'{ pfvf_port:1937  , pf:0 , vf:1937    , vf_active:1  },
'{ pfvf_port:1938  , pf:0 , vf:1938    , vf_active:1  },
'{ pfvf_port:1939  , pf:0 , vf:1939    , vf_active:1  },
'{ pfvf_port:1940  , pf:0 , vf:1940    , vf_active:1  },
'{ pfvf_port:1941  , pf:0 , vf:1941    , vf_active:1  },
'{ pfvf_port:1942  , pf:0 , vf:1942    , vf_active:1  },
'{ pfvf_port:1943  , pf:0 , vf:1943    , vf_active:1  },
'{ pfvf_port:1944  , pf:0 , vf:1944    , vf_active:1  },
'{ pfvf_port:1945  , pf:0 , vf:1945    , vf_active:1  },
'{ pfvf_port:1946  , pf:0 , vf:1946    , vf_active:1  },
'{ pfvf_port:1947  , pf:0 , vf:1947    , vf_active:1  },
'{ pfvf_port:1948  , pf:0 , vf:1948    , vf_active:1  },
'{ pfvf_port:1949  , pf:0 , vf:1949    , vf_active:1  },
'{ pfvf_port:1950  , pf:0 , vf:1950    , vf_active:1  },
'{ pfvf_port:1951  , pf:0 , vf:1951    , vf_active:1  },
'{ pfvf_port:1952  , pf:0 , vf:1952    , vf_active:1  },
'{ pfvf_port:1953  , pf:0 , vf:1953    , vf_active:1  },
'{ pfvf_port:1954  , pf:0 , vf:1954    , vf_active:1  },
'{ pfvf_port:1955  , pf:0 , vf:1955    , vf_active:1  },
'{ pfvf_port:1956  , pf:0 , vf:1956    , vf_active:1  },
'{ pfvf_port:1957  , pf:0 , vf:1957    , vf_active:1  },
'{ pfvf_port:1958  , pf:0 , vf:1958    , vf_active:1  },
'{ pfvf_port:1959  , pf:0 , vf:1959    , vf_active:1  },
'{ pfvf_port:1960  , pf:0 , vf:1960    , vf_active:1  },
'{ pfvf_port:1961  , pf:0 , vf:1961    , vf_active:1  },
'{ pfvf_port:1962  , pf:0 , vf:1962    , vf_active:1  },
'{ pfvf_port:1963  , pf:0 , vf:1963    , vf_active:1  },
'{ pfvf_port:1964  , pf:0 , vf:1964    , vf_active:1  },
'{ pfvf_port:1965  , pf:0 , vf:1965    , vf_active:1  },
'{ pfvf_port:1966  , pf:0 , vf:1966    , vf_active:1  },
'{ pfvf_port:1967  , pf:0 , vf:1967    , vf_active:1  },
'{ pfvf_port:1968  , pf:0 , vf:1968    , vf_active:1  },
'{ pfvf_port:1969  , pf:0 , vf:1969    , vf_active:1  },
'{ pfvf_port:1970  , pf:0 , vf:1970    , vf_active:1  },
'{ pfvf_port:1971  , pf:0 , vf:1971    , vf_active:1  },
'{ pfvf_port:1972  , pf:0 , vf:1972    , vf_active:1  },
'{ pfvf_port:1973  , pf:0 , vf:1973    , vf_active:1  },
'{ pfvf_port:1974  , pf:0 , vf:1974    , vf_active:1  },
'{ pfvf_port:1975  , pf:0 , vf:1975    , vf_active:1  },
'{ pfvf_port:1976  , pf:0 , vf:1976    , vf_active:1  },
'{ pfvf_port:1977  , pf:0 , vf:1977    , vf_active:1  },
'{ pfvf_port:1978  , pf:0 , vf:1978    , vf_active:1  },
'{ pfvf_port:1979  , pf:0 , vf:1979    , vf_active:1  },
'{ pfvf_port:1980  , pf:0 , vf:1980    , vf_active:1  },
'{ pfvf_port:1981  , pf:0 , vf:1981    , vf_active:1  },
'{ pfvf_port:1982  , pf:0 , vf:1982    , vf_active:1  },
'{ pfvf_port:1983  , pf:0 , vf:1983    , vf_active:1  },
'{ pfvf_port:1984  , pf:0 , vf:1984    , vf_active:1  },
'{ pfvf_port:1985  , pf:0 , vf:1985    , vf_active:1  },
'{ pfvf_port:1986  , pf:0 , vf:1986    , vf_active:1  },
'{ pfvf_port:1987  , pf:0 , vf:1987    , vf_active:1  },
'{ pfvf_port:1988  , pf:0 , vf:1988    , vf_active:1  },
'{ pfvf_port:1989  , pf:0 , vf:1989    , vf_active:1  },
'{ pfvf_port:1990  , pf:0 , vf:1990    , vf_active:1  },
'{ pfvf_port:1991  , pf:0 , vf:1991    , vf_active:1  },
'{ pfvf_port:1992  , pf:0 , vf:1992    , vf_active:1  },
'{ pfvf_port:1993  , pf:0 , vf:1993    , vf_active:1  },
'{ pfvf_port:1994  , pf:0 , vf:1994    , vf_active:1  },
'{ pfvf_port:1995  , pf:0 , vf:1995    , vf_active:1  },
'{ pfvf_port:1996  , pf:0 , vf:1996    , vf_active:1  },
'{ pfvf_port:1997  , pf:0 , vf:1997    , vf_active:1  },
'{ pfvf_port:1998  , pf:0 , vf:1998    , vf_active:1  },
'{ pfvf_port:1999  , pf:0 , vf:1999    , vf_active:1  },
'{ pfvf_port:2000  , pf:0 , vf:2000    , vf_active:1  },
'{ pfvf_port:2001  , pf:0 , vf:2001    , vf_active:1  },
'{ pfvf_port:2002  , pf:0 , vf:2002    , vf_active:1  },
'{ pfvf_port:2003  , pf:0 , vf:2003    , vf_active:1  },
'{ pfvf_port:2004  , pf:0 , vf:2004    , vf_active:1  },
'{ pfvf_port:2005  , pf:0 , vf:2005    , vf_active:1  },
'{ pfvf_port:2006  , pf:0 , vf:2006    , vf_active:1  },
'{ pfvf_port:2007  , pf:0 , vf:2007    , vf_active:1  },
'{ pfvf_port:2008  , pf:0 , vf:2008    , vf_active:1  },
'{ pfvf_port:2009  , pf:0 , vf:2009    , vf_active:1  },
'{ pfvf_port:2010  , pf:0 , vf:2010    , vf_active:1  },
'{ pfvf_port:2011  , pf:0 , vf:2011    , vf_active:1  },
'{ pfvf_port:2012  , pf:0 , vf:2012    , vf_active:1  },
'{ pfvf_port:2013  , pf:0 , vf:2013    , vf_active:1  },
'{ pfvf_port:2014  , pf:0 , vf:2014    , vf_active:1  },
'{ pfvf_port:2015  , pf:0 , vf:2015    , vf_active:1  },
'{ pfvf_port:2016  , pf:0 , vf:2016    , vf_active:1  },
'{ pfvf_port:2017  , pf:0 , vf:2017    , vf_active:1  },
'{ pfvf_port:2018  , pf:0 , vf:2018    , vf_active:1  },
'{ pfvf_port:2019  , pf:0 , vf:2019    , vf_active:1  },
'{ pfvf_port:2020  , pf:0 , vf:2020    , vf_active:1  },
'{ pfvf_port:2021  , pf:0 , vf:2021    , vf_active:1  },
'{ pfvf_port:2022  , pf:0 , vf:2022    , vf_active:1  },
'{ pfvf_port:2023  , pf:0 , vf:2023    , vf_active:1  },
'{ pfvf_port:2024  , pf:0 , vf:2024    , vf_active:1  },
'{ pfvf_port:2025  , pf:0 , vf:2025    , vf_active:1  },
'{ pfvf_port:2026  , pf:0 , vf:2026    , vf_active:1  },
'{ pfvf_port:2027  , pf:0 , vf:2027    , vf_active:1  },
'{ pfvf_port:2028  , pf:0 , vf:2028    , vf_active:1  },
'{ pfvf_port:2029  , pf:0 , vf:2029    , vf_active:1  },
'{ pfvf_port:2030  , pf:0 , vf:2030    , vf_active:1  },
'{ pfvf_port:2031  , pf:0 , vf:2031    , vf_active:1  },
'{ pfvf_port:2032  , pf:0 , vf:2032    , vf_active:1  },
'{ pfvf_port:2033  , pf:0 , vf:2033    , vf_active:1  },
'{ pfvf_port:2034  , pf:0 , vf:2034    , vf_active:1  },
'{ pfvf_port:2035  , pf:0 , vf:2035    , vf_active:1  },
'{ pfvf_port:2036  , pf:0 , vf:2036    , vf_active:1  },
'{ pfvf_port:2037  , pf:0 , vf:2037    , vf_active:1  },
'{ pfvf_port:2038  , pf:0 , vf:2038    , vf_active:1  },
'{ pfvf_port:2039  , pf:0 , vf:2039    , vf_active:1  },
'{ pfvf_port:2040  , pf:0 , vf:2040    , vf_active:1  },
'{ pfvf_port:2041  , pf:0 , vf:2041    , vf_active:1  },
'{ pfvf_port:2042  , pf:0 , vf:2042    , vf_active:1  },
'{ pfvf_port:2043  , pf:0 , vf:2043    , vf_active:1  },
'{ pfvf_port:2044  , pf:0 , vf:2044    , vf_active:1  },
'{ pfvf_port:2045  , pf:0 , vf:2045    , vf_active:1  },
'{ pfvf_port:2046  , pf:0 , vf:2046    , vf_active:1  },
'{ pfvf_port:2047  , pf:0 , vf:2047    , vf_active:1  }
        };
`endif


module top_tb;
  /** Parameter defines the clock frequency */
  parameter simulation_cycle = 50;

  //================================
  // Importing Required Packages 
  //================================
  import svt_axi_uvm_pkg::*;
  import uvm_pkg::*;
  
  //================================
  // Reset 
  //================================
  bit rst_n,clk;
  assign rst_n = axi_reset_if.reset;
  
	`ifdef DUMP
  initial 
  begin
    $vcdpluson;
    $vcdplusmemon();
  end
	`endif
  
  initial begin
     #1000;
     $display("TEST RUNNING\n");
  end
  
   /** Testbench 'System' Clock Generator */
  initial begin
    clk = 0 ;
    forever begin
      #(simulation_cycle/2)
        clk = ~clk ;
    end
  end

  //================================
  // VIP Interfaces
  //================================

  svt_axi_if axis_if_H();
  svt_axi_if axis_if_D();
  `ifndef TB_CONFIG_1
     `ifdef TB_CONFIG_4
       svt_axi_if TB4_axis_if_D0();
       svt_axi_if TB4_axis_if_D1();
       svt_axi_if TB4_axis_if_D2();
       svt_axi_if TB4_axis_if_D3();
    `else
      svt_axi_if axis_if_DN();
    `endif  
  `endif

  //================================
  // Coverage Interface
  //================================
  pf_vf_mux_if pf_vf_mux_cov_intf();

  /** TB Interface instance to provide access to the reset signal */
  axi_reset_if axi_reset_if();
  assign axi_reset_if.clk = clk;
  
  pcie_ss_axis_if #(
     .DATA_W (512),
     .USER_W (10)
  ) ho2mx_rx_remap (.clk(clk), .rst_n(rst_n));
  
  pcie_ss_axis_if #(
     .DATA_W (512),
     .USER_W (10)
  ) mx2ho_tx_remap(.clk(clk), .rst_n(rst_n));
   
  pcie_ss_axis_if #(
     .DATA_W (512),
     .USER_W (10)
  ) mx2fn_rx_remap[`NUM_PORT-1:0](.clk(clk), .rst_n(rst_n));
  
  pcie_ss_axis_if #(
     .DATA_W (512),
     .USER_W (10)
  ) fn2mx_tx_remap[`NUM_PORT-1:0](.clk(clk), .rst_n(rst_n));



	ofs_avst_if ofs_avst_if_inst();
  
  
  //================================
  // DUT Instantiation 
  //================================

  pf_vf_mux_w_params #(
     .MUX_NAME("A"),
     .NUM_RTABLE_ENTRIES(LOCAL_NUM_RTABLE_ENTRIES),
     .PFVF_ROUTING_TABLE(LOCAL_PFVF_ROUTING_TABLE)
  ) pf_vf_mux_a (
     .clk             (clk),
     .rst_n           (rst_n),
     .ho2mx_rx_port   (ho2mx_rx_remap),
     .mx2ho_tx_port   (mx2ho_tx_remap),
     .mx2fn_rx_port   (mx2fn_rx_remap),
     .fn2mx_tx_port   (fn2mx_tx_remap),
     .out_fifo_err    (),
     .out_fifo_perr   ()
  );
  
  `ifdef TB_CONFIG_1
    AXI_VIP AXI_VIP_INST(axis_if_D,axis_if_H);
  `elsif TB_CONFIG_4
    AXI_VIP AXI_VIP_INST(axis_if_D,axis_if_H,TB4_axis_if_D0,TB4_axis_if_D1,TB4_axis_if_D2,TB4_axis_if_D3);
  `else 
    AXI_VIP AXI_VIP_INST(axis_if_D,axis_if_DN,axis_if_H);
  `endif 
  
    initial begin
    /** Set the reset interface on the virtual sequencer */
    uvm_config_db#(virtual axi_reset_if.axi_reset_modport)::set(uvm_root::get(), "uvm_test_top.env.sequencer", "reset_mp", axi_reset_if.axi_reset_modport);
     uvm_config_db#(svt_axi_vif)::set(uvm_root::get(), "uvm_test_top.env.pf_vf_mux_system_env_H", "vif", axis_if_H);
     uvm_config_db#(svt_axi_vif)::set(uvm_root::get(), "uvm_test_top.env.pf_vf_mux_system_env_D", "vif", axis_if_D);
     `ifndef TB_CONFIG_1
        `ifdef TB_CONFIG_4
          uvm_config_db#(svt_axi_vif)::set(uvm_root::get(), "uvm_test_top.env.pf_vf_mux_system_env_TB4_D0", "vif", TB4_axis_if_D0);
          uvm_config_db#(svt_axi_vif)::set(uvm_root::get(), "uvm_test_top.env.pf_vf_mux_system_env_TB4_D1", "vif", TB4_axis_if_D1);
          uvm_config_db#(svt_axi_vif)::set(uvm_root::get(), "uvm_test_top.env.pf_vf_mux_system_env_TB4_D2", "vif", TB4_axis_if_D2);
          uvm_config_db#(svt_axi_vif)::set(uvm_root::get(), "uvm_test_top.env.pf_vf_mux_system_env_TB4_D3", "vif", TB4_axis_if_D3);
         `else 
          uvm_config_db#(svt_axi_vif)::set(uvm_root::get(), "uvm_test_top.env.pf_vf_mux_system_env_DN", "vif", axis_if_DN);
        `endif
     `endif  
     run_test();
     end

endmodule
