// Copyright 2022 Intel Corporation
// SPDX-License-Identifier: MIT

`include "ofs_plat_if.vh"

//
// Top level PIM-based module.
//

module ofs_plat_afu
   (
    // All platform wires, wrapped in one interface.
    ofs_plat_if plat_ifc
    );

    // ====================================================================
    //
    //  Get an AXI-MM host channel connection from the platform.
    //
    // ====================================================================

    // Up to two instances of HE LB will be created: one with EMIF and
    // one without.
`ifdef OFS_PLAT_PARAM_LOCAL_MEM_NUM_BANKS
    localparam NUM_ENG = (plat_ifc.host_chan.NUM_PORTS >= 2) ? 2 : 1;
`else
    // No local memory available
    localparam NUM_ENG = 1;
`endif

    // Instance of the PIM's standard AXI memory interface.
    ofs_plat_axi_mem_if
      #(
        // The PIM provides parameters for configuring a standard host
        // memory DMA AXI memory interface.
        `HOST_CHAN_AXI_MEM_PARAMS,
        // PIM interfaces can be configured to log traffic during
        // simulation. In ASE, see work/log_ofs_plat_host_chan.tsv.
        .LOG_CLASS(ofs_plat_log_pkg::HOST_CHAN)
        )
      axi_host_mem[NUM_ENG]();

    // Instance of the PIM's AXI memory lite interface, which will be
    // used to implement the AFU's CSR space.
    ofs_plat_axi_mem_lite_if
      #(
        // The AFU choses the data bus width of the interface and the
        // PIM adjusts the address space to match.
        `HOST_CHAN_AXI_MMIO_PARAMS(64),
        // Log MMIO traffic. (See the same parameter above on host_mem.)
        .LOG_CLASS(ofs_plat_log_pkg::HOST_CHAN)
        )
       axi_mmio64[NUM_ENG]();

    // HE LB's CSR interface is closer to Avalon, so the AXI-Lite CSR
    // interface is mapped to this.
    ofs_plat_avalon_mem_if
      #(
        `HOST_CHAN_AVALON_MMIO_PARAMS(64),
        .USER_WIDTH(axi_mmio64[0].USER_WIDTH + axi_mmio64[0].RID_WIDTH),
        .LOG_CLASS(ofs_plat_log_pkg::HOST_CHAN)
        )
      avmm_mmio64[NUM_ENG]();

    generate
        for (genvar p = 0; p < NUM_ENG; p = p + 1)
        begin : hc
            ofs_plat_host_chan_as_axi_mem_with_mmio
              #(
                // HE LB expects responses in order
                .SORT_READ_RESPONSES(1),
                .SORT_WRITE_RESPONSES(1)
                )
              primary_axi
               (
                .to_fiu(plat_ifc.host_chan.ports[p]),
                .host_mem_to_afu(axi_host_mem[p]),
                .mmio_to_afu(axi_mmio64[p]),

                .afu_clk(),
                .afu_reset_n()
                );

            // Map the AXI-Lite CSR interface to AVMM for use with the HE LB
            // CSR manager.
            assign avmm_mmio64[p].clk = axi_mmio64[p].clk;
            assign avmm_mmio64[p].reset_n = axi_mmio64[p].reset_n;
            assign avmm_mmio64[p].instance_number = axi_mmio64[p].instance_number;

            ofs_plat_axi_mem_lite_if_to_avalon_if
              #(
                // Clear the AXI user field in responses. It is unused,
                // so forcing it to 0 saves area.
                .PRESERVE_RESPONSE_USER(0),
                // Generate the AXI write response inside the shim.
                .LOCAL_WR_RESPONSE(1)
                )
              mmio_to_avmm
               (
                .axi_source(axi_mmio64[p]),
                .avmm_sink(avmm_mmio64[p])
                );

            // Tie off unused fields, including flow control. The HE LB CSR manager
            // is always ready and write responses are generated by the shim above.
            assign avmm_mmio64[p].waitrequest = 1'b0;
            assign avmm_mmio64[p].writeresponsevalid = 1'b0;
            assign avmm_mmio64[p].writeresponse = '0;
            assign avmm_mmio64[p].writeresponseuser = '0;
        end
    endgenerate


    // ====================================================================
    //
    //  Local memory
    //
    // ====================================================================

    // Two instances of ext_mem_if are defined. Only one will actually be
    // connected to a memory bank. The other is a dummy interface. This is
    // because two instances of he_lb_main() are instantiated. One will have
    // a local memory connection, the other will not.
    //
    // The HE_MEM_IDX macro, defined in filelist.txt, determines which
    // index has the real memory bank and which is the dummy.
    localparam HE_MEM_IDX = (`HE_MEM_IDX == 0) ? 0 : 1;
    localparam HE_LB_IDX = (HE_MEM_IDX == 0) ? 1 : 0;

`ifdef OFS_PLAT_PARAM_LOCAL_MEM_NUM_BANKS
    //
    // Local memory exists and the HE MEM instance has an available host port.
    //
    localparam HE_LB_EMIF_AVAIL = (HE_MEM_IDX < NUM_ENG);
    localparam HE_LB_EMIF_WIDTH = `OFS_PLAT_PARAM_LOCAL_MEM_DATA_WIDTH;

    // Local memory interface
    ofs_plat_axi_mem_if
      #(
        `LOCAL_MEM_AXI_MEM_PARAMS
        )
      ext_mem_if[NUM_ENG]();
`else
    //
    // No local memory
    //
    localparam HE_LB_EMIF_AVAIL = 0;
    localparam HE_LB_EMIF_WIDTH = 0;

    // Dummy memory interface, needed by he_lb_main.
    ofs_plat_axi_mem_if
      #(
        // Actual values here don't matter but some value is required
        .ADDR_WIDTH(10),
        .DATA_WIDTH(512)
        )
      ext_mem_if[NUM_ENG]();
`endif

    generate
        for (genvar p = 0; p < NUM_ENG; p = p + 1)
        begin : mem
            wire clk = axi_host_mem[p].clk;
            wire reset_n = axi_host_mem[p].reset_n;

            if ((p == HE_MEM_IDX) && (HE_LB_EMIF_AVAIL != 0))
            begin
                //
                // This engine is the HE MEM instance. Map bank 0 of local
                // memory to ext_mem_if[p].
                //
                ofs_plat_local_mem_as_axi_mem
                  #(
                    // Add a clock crossing
                    .ADD_CLOCK_CROSSING(1)
                    )
                  shim
                   (
                    .to_fiu(plat_ifc.local_mem.banks[0]),
                    .to_afu(ext_mem_if[p]),

                    .afu_clk(clk),
                    .afu_reset_n(reset_n)
                    );
            end
            else
            begin
                //
                // This engine is HE LB with no memory. Tie off the dummy
                // memory interface.
                //
                assign ext_mem_if[p].clk = clk;
                assign ext_mem_if[p].reset_n = reset_n;
                assign ext_mem_if[p].instance_number = 0;
                assign ext_mem_if[p].awready = 1'b1;
                assign ext_mem_if[p].wready = 1'b1;
                assign ext_mem_if[p].bvalid = 1'b0;
                assign ext_mem_if[p].arready = 1'b1;
                assign ext_mem_if[p].rvalid = 1'b0;
            end
        end
    endgenerate


    // ====================================================================
    //
    //  Tie off unused ports.
    //
    // ====================================================================

    // The PIM ties off unused devices, controlled by the AFU indicating
    // which devices it is using. This way, an AFU must know only about
    // the devices it uses. Tie-offs are thus portable, with the PIM
    // managing devices unused by and unknown to the AFU.
    ofs_plat_if_tie_off_unused
      #(
`ifdef OFS_PLAT_PARAM_LOCAL_MEM_NUM_BANKS
        // One bank of memory may be used
        .LOCAL_MEM_IN_USE_MASK(HE_LB_EMIF_AVAIL),
`endif
        // Up to 2 host channels are used, one for HE MEM and one for HE LB.
        // Turn the count into a bit mask.
        .HOST_CHAN_IN_USE_MASK((1 << NUM_ENG) - 1)
        )
        tie_off(plat_ifc);


    // =========================================================================
    //
    //   Instantiate the HE LB engines.
    //
    // =========================================================================

    generate
        for (genvar p = 0; p < NUM_ENG; p = p + 1)
        begin : eng
            wire clk = axi_host_mem[p].clk;
            wire reset_n = axi_host_mem[p].reset_n;

            // Connections to the CSR manager
            he_lb_pkg::he_csr_req  csr_req;
            he_lb_pkg::he_csr_dout csr_dout;
            he_lb_pkg::he_csr2eng  csr2eng;
            he_lb_pkg::he_eng2csr  eng2csr;

            // Use the PIM-generated AVMM interface for CSRs. AVMM
            // traffic will be merged into the host channel stream
            // by the PIM.

            assign csr_req.wen = avmm_mmio64[p].write;
            assign csr_req.ren = avmm_mmio64[p].read;
            // CSR manager addresses are to 32 bit chunks. The AVMM interface
            // addresses are to 64 bit chunks. For writes, if the first data byte
            // is unused then infer a 32 bit address in the high half of the 64
            // bit location. For reads, the HE LB CSR manager always expects
            // requests aligned to 64 bits.
            assign csr_req.addr = he_lb_pkg::CSR_AW'({ avmm_mmio64[p].address,
                                                       avmm_mmio64[p].write & ~avmm_mmio64[p].byteenable[0] });
            assign csr_req.din = avmm_mmio64[p].writedata;

            // Infer that a request is 64 bits when the first byte of
            // both 32 bit halves of a read or write or valid.
            assign csr_req.len = avmm_mmio64[p].byteenable[4] & avmm_mmio64[p].byteenable[0];

            assign csr_req.tag = he_lb_pkg::CSR_TAG_W'(avmm_mmio64[p].user);

            // Read responses from the CSR manager back to the AVMM interface
            assign avmm_mmio64[p].readdatavalid    = csr_dout.valid;    
            assign avmm_mmio64[p].readdata         = csr_dout.data;
            assign avmm_mmio64[p].response         = '0;
            assign avmm_mmio64[p].readresponseuser = csr_dout.tag;     


            // HE LB CSR manager
            he_lb_csr
              #(
                .CLK_MHZ(`OFS_PLAT_PARAM_CLOCKS_PCLK_FREQ),
                .HE_MEM_DATA_WIDTH((p == HE_MEM_IDX && HE_LB_EMIF_AVAIL != 0) ? HE_LB_EMIF_WIDTH : 0)
                )
              he_lb_csr
               (
                .clk,
                .rst_n(reset_n),

                .csr_req,
                .csr_dout,

                .csr2eng,
                .eng2csr
                );


            // Instantiate an HE LB engine
            he_lb_engines
              #(
                .EMIF(p == HE_MEM_IDX && HE_LB_EMIF_AVAIL != 0)
                )
              he_lb
               (
                .clk,
                .rst_n(reset_n),
                .csr2eng,
                .eng2csr,
                .axi_host_mem(axi_host_mem[p]),
                .emif_if(ext_mem_if[p])
                );
        end // block: eng
    endgenerate

endmodule
