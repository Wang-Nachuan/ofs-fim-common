// Copyright (C) 2023 Intel Corporation.
// SPDX-License-Identifier: MIT

//
// Description
//-----------------------------------------------------------------------------
//
// Common package for memory interface parameters. 
//
//-----------------------------------------------------------------------------

`ifndef __OFS_FIM_MEM_IF_PKG__
`define __OFS_FIM_MEM_IF_PKG__

// IP configuration database, generated by OFS script ofs_ip_cfg_db.tcl after
// IP generation.
`include "ofs_ip_cfg_db.vh"

package ofs_fim_mem_if_pkg;

   // FIM MEMORY PARAMS
   
   // Local memory interface bus width parameters:
   //
   // If no Memory Subsystem is present in the design or a type of memory interface isn't present in the subsystem component
   // then fallback values are selected for the parameters below.
   // The fallback values do not provide a functional mapping to IP interfaces. They are only defined for compilation
   // units included within common design files.

   // AXI-MM PARAMS
`ifdef OFS_FIM_IP_CFG_LOCAL_MEM_DEFINES_USER_AXI
   localparam NUM_MEM_CHANNELS        = `OFS_FIM_IP_CFG_LOCAL_MEM_NUM_AXI_CHANNELS;
   // AW
   parameter AXI_MEM_AWID_WIDTH       = `OFS_FIM_IP_CFG_LOCAL_MEM_AXI_AWID_WIDTH;
   parameter AXI_MEM_AWADDR_WIDTH     = `OFS_FIM_IP_CFG_LOCAL_MEM_AXI_AWADDR_WIDTH;
   parameter AXI_MEM_AWUSER_WIDTH     = `OFS_FIM_IP_CFG_LOCAL_MEM_AXI_AWUSER_WIDTH;
   // W
   parameter AXI_MEM_WDATA_WIDTH      = `OFS_FIM_IP_CFG_LOCAL_MEM_AXI_WDATA_WIDTH;
   parameter AXI_MEM_WUSER_WIDTH      = `OFS_FIM_IP_CFG_LOCAL_MEM_AXI_WUSER_WIDTH;
   // B
   parameter AXI_MEM_BID_WIDTH        = `OFS_FIM_IP_CFG_LOCAL_MEM_AXI_BID_WIDTH;
   parameter AXI_MEM_BUSER_WIDTH      = `OFS_FIM_IP_CFG_LOCAL_MEM_AXI_BUSER_WIDTH;
   // AR
   parameter AXI_MEM_ARID_WIDTH       = `OFS_FIM_IP_CFG_LOCAL_MEM_AXI_ARID_WIDTH;
   parameter AXI_MEM_ARADDR_WIDTH     = `OFS_FIM_IP_CFG_LOCAL_MEM_AXI_ARADDR_WIDTH;
   parameter AXI_MEM_ARUSER_WIDTH     = `OFS_FIM_IP_CFG_LOCAL_MEM_AXI_ARUSER_WIDTH;
   // R
   parameter AXI_MEM_RDATA_WIDTH      = `OFS_FIM_IP_CFG_LOCAL_MEM_AXI_RDATA_WIDTH;
   parameter AXI_MEM_RID_WIDTH        = `OFS_FIM_IP_CFG_LOCAL_MEM_AXI_RID_WIDTH;
   parameter AXI_MEM_RUSER_WIDTH      = `OFS_FIM_IP_CFG_LOCAL_MEM_AXI_RUSER_WIDTH;
`else 
   localparam NUM_MEM_CHANNELS        = 1;
   parameter AXI_MEM_AWID_WIDTH       = 1;
   parameter AXI_MEM_AWADDR_WIDTH     = 32;
   parameter AXI_MEM_AWUSER_WIDTH     = 1;
   parameter AXI_MEM_WDATA_WIDTH      = 512;
   parameter AXI_MEM_WUSER_WIDTH      = 1;
   parameter AXI_MEM_BID_WIDTH        = 1;
   parameter AXI_MEM_BUSER_WIDTH      = 1;
   parameter AXI_MEM_ARID_WIDTH       = 1;
   parameter AXI_MEM_ARADDR_WIDTH     = 32;
   parameter AXI_MEM_ARUSER_WIDTH     = 1;
   parameter AXI_MEM_RDATA_WIDTH      = 512;
   parameter AXI_MEM_RID_WIDTH        = 1;
   parameter AXI_MEM_RUSER_WIDTH      = 1;
`endif
   // This is defined by the AXI standard
   localparam AXI_MEM_BURST_LEN_WIDTH = 8;
   // TODO: Temporary
   localparam NUM_HBM_DEVICES = 2;

   // DDR4 PARAMS
`ifdef OFS_FIM_IP_CFG_LOCAL_MEM_DEFINES_EMIF_DDR4
   localparam NUM_DDR4_CHANNELS       = `OFS_FIM_IP_CFG_LOCAL_MEM_NUM_DDR4_CHANNELS;
   localparam DDR4_A_WIDTH            = `OFS_FIM_IP_CFG_LOCAL_MEM_DDR4_A_WIDTH;
   localparam DDR4_BA_WIDTH           = `OFS_FIM_IP_CFG_LOCAL_MEM_DDR4_BA_WIDTH;
   localparam DDR4_BG_WIDTH           = `OFS_FIM_IP_CFG_LOCAL_MEM_DDR4_BG_WIDTH;
   localparam DDR4_CK_WIDTH           = `OFS_FIM_IP_CFG_LOCAL_MEM_DDR4_CK_WIDTH;
   localparam DDR4_CKE_WIDTH          = `OFS_FIM_IP_CFG_LOCAL_MEM_DDR4_CKE_WIDTH;
   localparam DDR4_CS_WIDTH           = `OFS_FIM_IP_CFG_LOCAL_MEM_DDR4_CS_N_WIDTH;
   localparam DDR4_ODT_WIDTH          = `OFS_FIM_IP_CFG_LOCAL_MEM_DDR4_ODT_WIDTH;
   localparam DDR4_DQ_WIDTH           = `OFS_FIM_IP_CFG_LOCAL_MEM_DDR4_DQ_WIDTH;
`else
   localparam NUM_DDR4_CHANNELS       = 1;
   localparam DDR4_A_WIDTH            = 17;
   localparam DDR4_BA_WIDTH           = 2;
   localparam DDR4_BG_WIDTH           = 1;
   localparam DDR4_CK_WIDTH           = 1;
   localparam DDR4_CKE_WIDTH          = 1;
   localparam DDR4_CS_WIDTH           = 2;
   localparam DDR4_ODT_WIDTH          = 1;
   localparam DDR4_DQ_WIDTH           = 32;
`endif
   localparam DDR4_DQS_WIDTH          = DDR4_DQ_WIDTH/8;
   
`ifdef OFS_FIM_IP_CFG_LOCAL_MEM_DEFINES_HPS_DDR4
   localparam HPS_A_WIDTH            = `OFS_FIM_IP_CFG_LOCAL_MEM_HPS_A_WIDTH;
   localparam HPS_BA_WIDTH           = `OFS_FIM_IP_CFG_LOCAL_MEM_HPS_BA_WIDTH;
   localparam HPS_BG_WIDTH           = `OFS_FIM_IP_CFG_LOCAL_MEM_HPS_BG_WIDTH;
   localparam HPS_CK_WIDTH           = `OFS_FIM_IP_CFG_LOCAL_MEM_HPS_CK_WIDTH;
   localparam HPS_CKE_WIDTH          = `OFS_FIM_IP_CFG_LOCAL_MEM_HPS_CKE_WIDTH;
   localparam HPS_CS_WIDTH           = `OFS_FIM_IP_CFG_LOCAL_MEM_HPS_CS_N_WIDTH;
   localparam HPS_ODT_WIDTH          = `OFS_FIM_IP_CFG_LOCAL_MEM_HPS_ODT_WIDTH;
   localparam HPS_DQ_WIDTH           = `OFS_FIM_IP_CFG_LOCAL_MEM_HPS_DQ_WIDTH;
`else
   localparam NUM_HPS_CHANNELS       = 1;
   localparam HPS_A_WIDTH            = 17;
   localparam HPS_BA_WIDTH           = 2;
   localparam HPS_BG_WIDTH           = 1;
   localparam HPS_CK_WIDTH           = 1;
   localparam HPS_CKE_WIDTH          = 1;
   localparam HPS_CS_WIDTH           = 2;
   localparam HPS_ODT_WIDTH          = 1;
   localparam HPS_DQ_WIDTH           = 32;
`endif
   localparam HPS_DQS_WIDTH          = HPS_DQ_WIDTH/8;
   
endpackage : ofs_fim_mem_if_pkg

`endif //  `ifndef __OFS_FIM_MEM_IF_PKG__
   
